magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 16 21 1159 203
rect 29 -17 63 21
<< scnmos >>
rect 103 47 133 177
rect 187 47 217 177
rect 271 47 301 177
rect 355 47 385 177
rect 439 47 469 177
rect 627 47 657 177
rect 711 47 741 177
rect 795 47 825 177
rect 879 47 909 177
rect 963 47 993 177
rect 1047 47 1077 177
<< scpmoshvt >>
rect 103 297 133 497
rect 187 297 217 497
rect 271 297 301 497
rect 355 297 385 497
rect 439 297 469 497
rect 523 297 553 497
rect 607 297 637 497
rect 795 297 825 497
rect 879 297 909 497
rect 963 297 993 497
rect 1047 297 1077 497
<< ndiff >>
rect 42 163 103 177
rect 42 129 59 163
rect 93 129 103 163
rect 42 95 103 129
rect 42 61 59 95
rect 93 61 103 95
rect 42 47 103 61
rect 133 163 187 177
rect 133 129 143 163
rect 177 129 187 163
rect 133 95 187 129
rect 133 61 143 95
rect 177 61 187 95
rect 133 47 187 61
rect 217 163 271 177
rect 217 129 227 163
rect 261 129 271 163
rect 217 95 271 129
rect 217 61 227 95
rect 261 61 271 95
rect 217 47 271 61
rect 301 95 355 177
rect 301 61 311 95
rect 345 61 355 95
rect 301 47 355 61
rect 385 163 439 177
rect 385 129 395 163
rect 429 129 439 163
rect 385 95 439 129
rect 385 61 395 95
rect 429 61 439 95
rect 385 47 439 61
rect 469 95 521 177
rect 469 61 479 95
rect 513 61 521 95
rect 469 47 521 61
rect 575 95 627 177
rect 575 61 583 95
rect 617 61 627 95
rect 575 47 627 61
rect 657 163 711 177
rect 657 129 667 163
rect 701 129 711 163
rect 657 47 711 129
rect 741 163 795 177
rect 741 129 751 163
rect 785 129 795 163
rect 741 95 795 129
rect 741 61 751 95
rect 785 61 795 95
rect 741 47 795 61
rect 825 95 879 177
rect 825 61 835 95
rect 869 61 879 95
rect 825 47 879 61
rect 909 163 963 177
rect 909 129 919 163
rect 953 129 963 163
rect 909 95 963 129
rect 909 61 919 95
rect 953 61 963 95
rect 909 47 963 61
rect 993 95 1047 177
rect 993 61 1003 95
rect 1037 61 1047 95
rect 993 47 1047 61
rect 1077 163 1133 177
rect 1077 129 1087 163
rect 1121 129 1133 163
rect 1077 95 1133 129
rect 1077 61 1087 95
rect 1121 61 1133 95
rect 1077 47 1133 61
<< pdiff >>
rect 27 477 103 497
rect 27 443 53 477
rect 87 443 103 477
rect 27 409 103 443
rect 27 375 53 409
rect 87 375 103 409
rect 27 341 103 375
rect 27 307 53 341
rect 87 307 103 341
rect 27 297 103 307
rect 133 477 187 497
rect 133 443 143 477
rect 177 443 187 477
rect 133 297 187 443
rect 217 341 271 497
rect 217 307 227 341
rect 261 307 271 341
rect 217 297 271 307
rect 301 477 355 497
rect 301 443 311 477
rect 345 443 355 477
rect 301 297 355 443
rect 385 341 439 497
rect 385 307 395 341
rect 429 307 439 341
rect 385 297 439 307
rect 469 477 523 497
rect 469 443 479 477
rect 513 443 523 477
rect 469 297 523 443
rect 553 477 607 497
rect 553 443 563 477
rect 597 443 607 477
rect 553 409 607 443
rect 553 375 563 409
rect 597 375 607 409
rect 553 297 607 375
rect 637 477 689 497
rect 637 443 647 477
rect 681 443 689 477
rect 637 297 689 443
rect 743 477 795 497
rect 743 443 751 477
rect 785 443 795 477
rect 743 297 795 443
rect 825 409 879 497
rect 825 375 835 409
rect 869 375 879 409
rect 825 341 879 375
rect 825 307 835 341
rect 869 307 879 341
rect 825 297 879 307
rect 909 477 963 497
rect 909 443 919 477
rect 953 443 963 477
rect 909 409 963 443
rect 909 375 919 409
rect 953 375 963 409
rect 909 341 963 375
rect 909 307 919 341
rect 953 307 963 341
rect 909 297 963 307
rect 993 485 1047 497
rect 993 451 1003 485
rect 1037 451 1047 485
rect 993 417 1047 451
rect 993 383 1003 417
rect 1037 383 1047 417
rect 993 297 1047 383
rect 1077 477 1133 497
rect 1077 443 1087 477
rect 1121 443 1133 477
rect 1077 409 1133 443
rect 1077 375 1087 409
rect 1121 375 1133 409
rect 1077 341 1133 375
rect 1077 307 1087 341
rect 1121 307 1133 341
rect 1077 297 1133 307
<< ndiffc >>
rect 59 129 93 163
rect 59 61 93 95
rect 143 129 177 163
rect 143 61 177 95
rect 227 129 261 163
rect 227 61 261 95
rect 311 61 345 95
rect 395 129 429 163
rect 395 61 429 95
rect 479 61 513 95
rect 583 61 617 95
rect 667 129 701 163
rect 751 129 785 163
rect 751 61 785 95
rect 835 61 869 95
rect 919 129 953 163
rect 919 61 953 95
rect 1003 61 1037 95
rect 1087 129 1121 163
rect 1087 61 1121 95
<< pdiffc >>
rect 53 443 87 477
rect 53 375 87 409
rect 53 307 87 341
rect 143 443 177 477
rect 227 307 261 341
rect 311 443 345 477
rect 395 307 429 341
rect 479 443 513 477
rect 563 443 597 477
rect 563 375 597 409
rect 647 443 681 477
rect 751 443 785 477
rect 835 375 869 409
rect 835 307 869 341
rect 919 443 953 477
rect 919 375 953 409
rect 919 307 953 341
rect 1003 451 1037 485
rect 1003 383 1037 417
rect 1087 443 1121 477
rect 1087 375 1121 409
rect 1087 307 1121 341
<< poly >>
rect 103 497 133 523
rect 187 497 217 523
rect 271 497 301 523
rect 355 497 385 523
rect 439 497 469 523
rect 523 497 553 523
rect 607 497 637 523
rect 795 497 825 523
rect 879 497 909 523
rect 963 497 993 523
rect 1047 497 1077 523
rect 103 265 133 297
rect 187 265 217 297
rect 271 265 301 297
rect 355 265 385 297
rect 439 265 469 297
rect 91 249 145 265
rect 91 215 101 249
rect 135 215 145 249
rect 91 199 145 215
rect 187 249 469 265
rect 187 215 343 249
rect 377 215 411 249
rect 445 215 469 249
rect 187 199 469 215
rect 523 265 553 297
rect 607 265 637 297
rect 795 265 825 297
rect 879 265 909 297
rect 523 249 741 265
rect 523 215 577 249
rect 611 215 741 249
rect 523 199 741 215
rect 103 177 133 199
rect 187 177 217 199
rect 271 177 301 199
rect 355 177 385 199
rect 439 177 469 199
rect 627 177 657 199
rect 711 177 741 199
rect 795 249 909 265
rect 795 215 835 249
rect 869 215 909 249
rect 795 199 909 215
rect 795 177 825 199
rect 879 177 909 199
rect 963 265 993 297
rect 1047 265 1077 297
rect 963 249 1077 265
rect 963 215 1014 249
rect 1048 215 1077 249
rect 963 199 1077 215
rect 963 177 993 199
rect 1047 177 1077 199
rect 103 21 133 47
rect 187 21 217 47
rect 271 21 301 47
rect 355 21 385 47
rect 439 21 469 47
rect 627 21 657 47
rect 711 21 741 47
rect 795 21 825 47
rect 879 21 909 47
rect 963 21 993 47
rect 1047 21 1077 47
<< polycont >>
rect 101 215 135 249
rect 343 215 377 249
rect 411 215 445 249
rect 577 215 611 249
rect 835 215 869 249
rect 1014 215 1048 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 477 87 493
rect 17 443 53 477
rect 127 477 193 527
rect 127 443 143 477
rect 177 443 193 477
rect 295 477 361 527
rect 295 443 311 477
rect 345 443 361 477
rect 463 477 529 527
rect 463 443 479 477
rect 513 443 529 477
rect 563 477 597 493
rect 17 409 87 443
rect 563 409 597 443
rect 640 477 690 527
rect 640 443 647 477
rect 681 443 690 477
rect 640 427 690 443
rect 737 477 953 493
rect 737 443 751 477
rect 785 459 919 477
rect 737 427 785 443
rect 17 375 53 409
rect 87 375 513 409
rect 17 341 87 375
rect 17 307 53 341
rect 17 291 87 307
rect 17 171 51 291
rect 121 257 177 341
rect 85 249 177 257
rect 85 215 101 249
rect 135 215 177 249
rect 211 307 227 341
rect 261 307 395 341
rect 429 307 445 341
rect 211 289 445 307
rect 479 323 513 375
rect 827 409 876 425
rect 827 393 835 409
rect 597 375 835 393
rect 869 375 876 409
rect 563 359 876 375
rect 479 289 581 323
rect 211 181 291 289
rect 325 249 513 255
rect 325 215 343 249
rect 377 215 411 249
rect 445 215 513 249
rect 547 249 581 289
rect 547 215 577 249
rect 611 215 627 249
rect 17 163 109 171
rect 17 129 59 163
rect 93 129 109 163
rect 17 95 109 129
rect 17 61 59 95
rect 93 61 109 95
rect 17 53 109 61
rect 143 163 177 181
rect 143 95 177 129
rect 143 17 177 61
rect 211 163 445 181
rect 211 129 227 163
rect 261 145 395 163
rect 261 129 277 145
rect 211 95 277 129
rect 379 129 395 145
rect 429 129 445 163
rect 479 179 513 215
rect 679 179 717 359
rect 827 341 876 359
rect 827 307 835 341
rect 869 307 876 341
rect 827 289 876 307
rect 919 409 953 443
rect 919 341 953 375
rect 987 485 1053 527
rect 987 451 1003 485
rect 1037 451 1053 485
rect 987 417 1053 451
rect 987 383 1003 417
rect 1037 383 1053 417
rect 987 367 1053 383
rect 1087 477 1142 493
rect 1121 443 1142 477
rect 1087 409 1142 443
rect 1121 375 1142 409
rect 1087 341 1142 375
rect 953 307 1087 333
rect 1121 307 1142 341
rect 919 291 1142 307
rect 756 249 964 255
rect 756 215 835 249
rect 869 215 964 249
rect 998 249 1179 255
rect 998 215 1014 249
rect 1048 215 1179 249
rect 479 163 717 179
rect 479 145 667 163
rect 647 129 667 145
rect 701 129 717 163
rect 751 163 1142 181
rect 785 145 919 163
rect 785 129 801 145
rect 211 61 227 95
rect 261 61 277 95
rect 211 51 277 61
rect 311 95 345 111
rect 311 17 345 61
rect 379 95 445 129
rect 379 61 395 95
rect 429 61 445 95
rect 379 51 445 61
rect 479 95 513 111
rect 751 95 801 129
rect 903 129 919 145
rect 953 145 1087 163
rect 953 129 969 145
rect 479 17 513 61
rect 561 61 583 95
rect 617 61 751 95
rect 785 61 801 95
rect 561 51 801 61
rect 835 95 869 111
rect 835 17 869 61
rect 903 95 969 129
rect 1071 129 1087 145
rect 1121 129 1142 163
rect 903 61 919 95
rect 953 61 969 95
rect 903 51 969 61
rect 1003 95 1037 111
rect 1003 17 1037 61
rect 1071 95 1142 129
rect 1071 61 1087 95
rect 1121 61 1142 95
rect 1071 53 1142 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 121 221 155 255 0 FreeSans 400 180 0 0 B1_N
port 3 nsew signal input
flabel locali s 1041 221 1075 255 0 FreeSans 400 180 0 0 A1
port 1 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 400 180 0 0 A2
port 2 nsew signal input
flabel locali s 397 85 431 119 0 FreeSans 400 180 0 0 X
port 8 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o21ba_4
rlabel metal1 s 0 -48 1196 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 1328502
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1319502
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 5.980 0.000 
<< end >>
