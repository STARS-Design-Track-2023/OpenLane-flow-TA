magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 696 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 267 47 297 177
rect 362 47 392 177
rect 480 47 510 177
rect 580 47 610 177
<< scpmoshvt >>
rect 79 297 109 497
rect 267 297 297 497
rect 362 297 392 497
rect 480 297 510 497
rect 580 297 610 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 161 161 177
rect 109 127 119 161
rect 153 127 161 161
rect 109 93 161 127
rect 109 59 119 93
rect 153 59 161 93
rect 109 47 161 59
rect 215 161 267 177
rect 215 127 223 161
rect 257 127 267 161
rect 215 93 267 127
rect 215 59 223 93
rect 257 59 267 93
rect 215 47 267 59
rect 297 93 362 177
rect 297 59 313 93
rect 347 59 362 93
rect 297 47 362 59
rect 392 161 480 177
rect 392 127 402 161
rect 436 127 480 161
rect 392 93 480 127
rect 392 59 402 93
rect 436 59 480 93
rect 392 47 480 59
rect 510 47 580 177
rect 610 161 670 177
rect 610 127 628 161
rect 662 127 670 161
rect 610 93 670 127
rect 610 59 628 93
rect 662 59 670 93
rect 610 47 670 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 161 497
rect 109 451 119 485
rect 153 451 161 485
rect 109 417 161 451
rect 109 383 119 417
rect 153 383 161 417
rect 109 349 161 383
rect 109 315 119 349
rect 153 315 161 349
rect 109 297 161 315
rect 215 485 267 497
rect 215 451 223 485
rect 257 451 267 485
rect 215 417 267 451
rect 215 383 223 417
rect 257 383 267 417
rect 215 297 267 383
rect 297 297 362 497
rect 392 485 480 497
rect 392 451 402 485
rect 436 451 480 485
rect 392 417 480 451
rect 392 383 402 417
rect 436 383 480 417
rect 392 349 480 383
rect 392 315 402 349
rect 436 315 480 349
rect 392 297 480 315
rect 510 485 580 497
rect 510 451 528 485
rect 562 451 580 485
rect 510 417 580 451
rect 510 383 528 417
rect 562 383 580 417
rect 510 297 580 383
rect 610 485 670 497
rect 610 451 628 485
rect 662 451 670 485
rect 610 417 670 451
rect 610 383 628 417
rect 662 383 670 417
rect 610 349 670 383
rect 610 315 628 349
rect 662 315 670 349
rect 610 297 670 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 127 153 161
rect 119 59 153 93
rect 223 127 257 161
rect 223 59 257 93
rect 313 59 347 93
rect 402 127 436 161
rect 402 59 436 93
rect 628 127 662 161
rect 628 59 662 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 223 451 257 485
rect 223 383 257 417
rect 402 451 436 485
rect 402 383 436 417
rect 402 315 436 349
rect 528 451 562 485
rect 528 383 562 417
rect 628 451 662 485
rect 628 383 662 417
rect 628 315 662 349
<< poly >>
rect 79 497 109 523
rect 267 497 297 523
rect 362 497 392 523
rect 480 497 510 523
rect 580 497 610 523
rect 79 259 109 297
rect 267 265 297 297
rect 362 265 392 297
rect 480 265 510 297
rect 580 265 610 297
rect 79 249 152 259
rect 79 215 102 249
rect 136 215 152 249
rect 79 205 152 215
rect 266 249 320 265
rect 266 215 276 249
rect 310 215 320 249
rect 79 177 109 205
rect 266 199 320 215
rect 362 249 438 265
rect 362 215 394 249
rect 428 215 438 249
rect 362 199 438 215
rect 480 249 538 265
rect 480 215 494 249
rect 528 215 538 249
rect 480 199 538 215
rect 580 249 715 265
rect 580 215 665 249
rect 699 215 715 249
rect 580 199 715 215
rect 267 177 297 199
rect 362 177 392 199
rect 480 177 510 199
rect 580 177 610 199
rect 79 21 109 47
rect 267 21 297 47
rect 362 21 392 47
rect 480 21 510 47
rect 580 21 610 47
<< polycont >>
rect 102 215 136 249
rect 276 215 310 249
rect 394 215 428 249
rect 494 215 528 249
rect 665 215 699 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 485 85 493
rect 17 451 35 485
rect 69 451 85 485
rect 17 417 85 451
rect 17 383 35 417
rect 69 383 85 417
rect 17 349 85 383
rect 17 315 35 349
rect 69 315 85 349
rect 17 299 85 315
rect 119 485 153 527
rect 119 417 153 451
rect 119 349 153 383
rect 207 485 257 527
rect 207 451 223 485
rect 207 417 257 451
rect 207 383 223 417
rect 207 367 257 383
rect 386 485 452 493
rect 386 451 402 485
rect 436 451 452 485
rect 386 417 452 451
rect 386 383 402 417
rect 436 383 452 417
rect 386 349 452 383
rect 512 485 578 527
rect 512 451 528 485
rect 562 451 578 485
rect 512 417 578 451
rect 512 383 528 417
rect 562 383 578 417
rect 512 367 578 383
rect 612 485 678 493
rect 612 451 628 485
rect 662 451 678 485
rect 612 417 678 451
rect 612 383 628 417
rect 662 383 678 417
rect 386 333 402 349
rect 119 299 153 315
rect 191 315 402 333
rect 436 333 452 349
rect 612 349 678 383
rect 612 333 628 349
rect 436 315 628 333
rect 662 315 678 349
rect 191 299 678 315
rect 17 177 52 299
rect 191 249 225 299
rect 86 215 102 249
rect 136 215 225 249
rect 260 249 344 255
rect 260 215 276 249
rect 310 215 344 249
rect 378 249 444 255
rect 378 215 394 249
rect 428 215 444 249
rect 478 249 544 255
rect 478 215 494 249
rect 528 215 544 249
rect 17 161 85 177
rect 17 127 35 161
rect 69 127 85 161
rect 17 93 85 127
rect 17 59 35 93
rect 69 59 85 93
rect 17 51 85 59
rect 119 161 169 177
rect 153 127 169 161
rect 119 93 169 127
rect 153 59 169 93
rect 119 17 169 59
rect 207 161 452 181
rect 207 127 223 161
rect 257 147 402 161
rect 257 127 273 147
rect 207 93 273 127
rect 386 127 402 147
rect 436 127 452 161
rect 207 59 223 93
rect 257 59 273 93
rect 207 51 273 59
rect 307 93 352 109
rect 307 59 313 93
rect 347 59 352 93
rect 307 17 352 59
rect 386 93 452 127
rect 386 59 402 93
rect 436 59 452 93
rect 386 51 452 59
rect 578 173 612 299
rect 649 249 719 265
rect 649 215 665 249
rect 699 215 719 249
rect 578 161 678 173
rect 578 127 628 161
rect 662 127 678 161
rect 578 93 678 127
rect 578 59 628 93
rect 662 59 678 93
rect 578 51 678 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 673 221 707 255 0 FreeSans 250 0 0 0 C1
port 4 nsew signal input
flabel locali s 494 221 528 255 0 FreeSans 250 0 0 0 B1
port 3 nsew signal input
flabel locali s 402 221 436 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 310 221 344 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 30 85 64 119 0 FreeSans 250 0 0 0 X
port 9 nsew signal output
flabel locali s 30 425 64 459 0 FreeSans 250 0 0 0 X
port 9 nsew signal output
flabel locali s 30 357 64 391 0 FreeSans 250 0 0 0 X
port 9 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o211a_1
rlabel metal1 s 0 -48 736 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 755464
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 748680
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.680 0.000 
<< end >>
