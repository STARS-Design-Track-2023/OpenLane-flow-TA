magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< pwell >>
rect 15 163 811 1225
<< nmoslvt >>
rect 171 189 201 1199
rect 257 189 293 1199
rect 349 189 385 1199
rect 441 189 477 1199
rect 533 189 569 1199
rect 625 189 655 1199
<< ndiff >>
rect 111 1187 171 1199
rect 111 1153 126 1187
rect 160 1153 171 1187
rect 111 1119 171 1153
rect 111 1085 126 1119
rect 160 1085 171 1119
rect 111 1051 171 1085
rect 111 1017 126 1051
rect 160 1017 171 1051
rect 111 983 171 1017
rect 111 949 126 983
rect 160 949 171 983
rect 111 915 171 949
rect 111 881 126 915
rect 160 881 171 915
rect 111 847 171 881
rect 111 813 126 847
rect 160 813 171 847
rect 111 779 171 813
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 1187 257 1199
rect 201 1153 212 1187
rect 246 1153 257 1187
rect 201 1119 257 1153
rect 201 1085 212 1119
rect 246 1085 257 1119
rect 201 1051 257 1085
rect 201 1017 212 1051
rect 246 1017 257 1051
rect 201 983 257 1017
rect 201 949 212 983
rect 246 949 257 983
rect 201 915 257 949
rect 201 881 212 915
rect 246 881 257 915
rect 201 847 257 881
rect 201 813 212 847
rect 246 813 257 847
rect 201 779 257 813
rect 201 745 212 779
rect 246 745 257 779
rect 201 711 257 745
rect 201 677 212 711
rect 246 677 257 711
rect 201 643 257 677
rect 201 609 212 643
rect 246 609 257 643
rect 201 575 257 609
rect 201 541 212 575
rect 246 541 257 575
rect 201 507 257 541
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 293 1187 349 1199
rect 293 1153 304 1187
rect 338 1153 349 1187
rect 293 1119 349 1153
rect 293 1085 304 1119
rect 338 1085 349 1119
rect 293 1051 349 1085
rect 293 1017 304 1051
rect 338 1017 349 1051
rect 293 983 349 1017
rect 293 949 304 983
rect 338 949 349 983
rect 293 915 349 949
rect 293 881 304 915
rect 338 881 349 915
rect 293 847 349 881
rect 293 813 304 847
rect 338 813 349 847
rect 293 779 349 813
rect 293 745 304 779
rect 338 745 349 779
rect 293 711 349 745
rect 293 677 304 711
rect 338 677 349 711
rect 293 643 349 677
rect 293 609 304 643
rect 338 609 349 643
rect 293 575 349 609
rect 293 541 304 575
rect 338 541 349 575
rect 293 507 349 541
rect 293 473 304 507
rect 338 473 349 507
rect 293 439 349 473
rect 293 405 304 439
rect 338 405 349 439
rect 293 371 349 405
rect 293 337 304 371
rect 338 337 349 371
rect 293 303 349 337
rect 293 269 304 303
rect 338 269 349 303
rect 293 235 349 269
rect 293 201 304 235
rect 338 201 349 235
rect 293 189 349 201
rect 385 1187 441 1199
rect 385 1153 396 1187
rect 430 1153 441 1187
rect 385 1119 441 1153
rect 385 1085 396 1119
rect 430 1085 441 1119
rect 385 1051 441 1085
rect 385 1017 396 1051
rect 430 1017 441 1051
rect 385 983 441 1017
rect 385 949 396 983
rect 430 949 441 983
rect 385 915 441 949
rect 385 881 396 915
rect 430 881 441 915
rect 385 847 441 881
rect 385 813 396 847
rect 430 813 441 847
rect 385 779 441 813
rect 385 745 396 779
rect 430 745 441 779
rect 385 711 441 745
rect 385 677 396 711
rect 430 677 441 711
rect 385 643 441 677
rect 385 609 396 643
rect 430 609 441 643
rect 385 575 441 609
rect 385 541 396 575
rect 430 541 441 575
rect 385 507 441 541
rect 385 473 396 507
rect 430 473 441 507
rect 385 439 441 473
rect 385 405 396 439
rect 430 405 441 439
rect 385 371 441 405
rect 385 337 396 371
rect 430 337 441 371
rect 385 303 441 337
rect 385 269 396 303
rect 430 269 441 303
rect 385 235 441 269
rect 385 201 396 235
rect 430 201 441 235
rect 385 189 441 201
rect 477 1187 533 1199
rect 477 1153 488 1187
rect 522 1153 533 1187
rect 477 1119 533 1153
rect 477 1085 488 1119
rect 522 1085 533 1119
rect 477 1051 533 1085
rect 477 1017 488 1051
rect 522 1017 533 1051
rect 477 983 533 1017
rect 477 949 488 983
rect 522 949 533 983
rect 477 915 533 949
rect 477 881 488 915
rect 522 881 533 915
rect 477 847 533 881
rect 477 813 488 847
rect 522 813 533 847
rect 477 779 533 813
rect 477 745 488 779
rect 522 745 533 779
rect 477 711 533 745
rect 477 677 488 711
rect 522 677 533 711
rect 477 643 533 677
rect 477 609 488 643
rect 522 609 533 643
rect 477 575 533 609
rect 477 541 488 575
rect 522 541 533 575
rect 477 507 533 541
rect 477 473 488 507
rect 522 473 533 507
rect 477 439 533 473
rect 477 405 488 439
rect 522 405 533 439
rect 477 371 533 405
rect 477 337 488 371
rect 522 337 533 371
rect 477 303 533 337
rect 477 269 488 303
rect 522 269 533 303
rect 477 235 533 269
rect 477 201 488 235
rect 522 201 533 235
rect 477 189 533 201
rect 569 1187 625 1199
rect 569 1153 580 1187
rect 614 1153 625 1187
rect 569 1119 625 1153
rect 569 1085 580 1119
rect 614 1085 625 1119
rect 569 1051 625 1085
rect 569 1017 580 1051
rect 614 1017 625 1051
rect 569 983 625 1017
rect 569 949 580 983
rect 614 949 625 983
rect 569 915 625 949
rect 569 881 580 915
rect 614 881 625 915
rect 569 847 625 881
rect 569 813 580 847
rect 614 813 625 847
rect 569 779 625 813
rect 569 745 580 779
rect 614 745 625 779
rect 569 711 625 745
rect 569 677 580 711
rect 614 677 625 711
rect 569 643 625 677
rect 569 609 580 643
rect 614 609 625 643
rect 569 575 625 609
rect 569 541 580 575
rect 614 541 625 575
rect 569 507 625 541
rect 569 473 580 507
rect 614 473 625 507
rect 569 439 625 473
rect 569 405 580 439
rect 614 405 625 439
rect 569 371 625 405
rect 569 337 580 371
rect 614 337 625 371
rect 569 303 625 337
rect 569 269 580 303
rect 614 269 625 303
rect 569 235 625 269
rect 569 201 580 235
rect 614 201 625 235
rect 569 189 625 201
rect 655 1187 715 1199
rect 655 1153 666 1187
rect 700 1153 715 1187
rect 655 1119 715 1153
rect 655 1085 666 1119
rect 700 1085 715 1119
rect 655 1051 715 1085
rect 655 1017 666 1051
rect 700 1017 715 1051
rect 655 983 715 1017
rect 655 949 666 983
rect 700 949 715 983
rect 655 915 715 949
rect 655 881 666 915
rect 700 881 715 915
rect 655 847 715 881
rect 655 813 666 847
rect 700 813 715 847
rect 655 779 715 813
rect 655 745 666 779
rect 700 745 715 779
rect 655 711 715 745
rect 655 677 666 711
rect 700 677 715 711
rect 655 643 715 677
rect 655 609 666 643
rect 700 609 715 643
rect 655 575 715 609
rect 655 541 666 575
rect 700 541 715 575
rect 655 507 715 541
rect 655 473 666 507
rect 700 473 715 507
rect 655 439 715 473
rect 655 405 666 439
rect 700 405 715 439
rect 655 371 715 405
rect 655 337 666 371
rect 700 337 715 371
rect 655 303 715 337
rect 655 269 666 303
rect 700 269 715 303
rect 655 235 715 269
rect 655 201 666 235
rect 700 201 715 235
rect 655 189 715 201
<< ndiffc >>
rect 126 1153 160 1187
rect 126 1085 160 1119
rect 126 1017 160 1051
rect 126 949 160 983
rect 126 881 160 915
rect 126 813 160 847
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 1153 246 1187
rect 212 1085 246 1119
rect 212 1017 246 1051
rect 212 949 246 983
rect 212 881 246 915
rect 212 813 246 847
rect 212 745 246 779
rect 212 677 246 711
rect 212 609 246 643
rect 212 541 246 575
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 304 1153 338 1187
rect 304 1085 338 1119
rect 304 1017 338 1051
rect 304 949 338 983
rect 304 881 338 915
rect 304 813 338 847
rect 304 745 338 779
rect 304 677 338 711
rect 304 609 338 643
rect 304 541 338 575
rect 304 473 338 507
rect 304 405 338 439
rect 304 337 338 371
rect 304 269 338 303
rect 304 201 338 235
rect 396 1153 430 1187
rect 396 1085 430 1119
rect 396 1017 430 1051
rect 396 949 430 983
rect 396 881 430 915
rect 396 813 430 847
rect 396 745 430 779
rect 396 677 430 711
rect 396 609 430 643
rect 396 541 430 575
rect 396 473 430 507
rect 396 405 430 439
rect 396 337 430 371
rect 396 269 430 303
rect 396 201 430 235
rect 488 1153 522 1187
rect 488 1085 522 1119
rect 488 1017 522 1051
rect 488 949 522 983
rect 488 881 522 915
rect 488 813 522 847
rect 488 745 522 779
rect 488 677 522 711
rect 488 609 522 643
rect 488 541 522 575
rect 488 473 522 507
rect 488 405 522 439
rect 488 337 522 371
rect 488 269 522 303
rect 488 201 522 235
rect 580 1153 614 1187
rect 580 1085 614 1119
rect 580 1017 614 1051
rect 580 949 614 983
rect 580 881 614 915
rect 580 813 614 847
rect 580 745 614 779
rect 580 677 614 711
rect 580 609 614 643
rect 580 541 614 575
rect 580 473 614 507
rect 580 405 614 439
rect 580 337 614 371
rect 580 269 614 303
rect 580 201 614 235
rect 666 1153 700 1187
rect 666 1085 700 1119
rect 666 1017 700 1051
rect 666 949 700 983
rect 666 881 700 915
rect 666 813 700 847
rect 666 745 700 779
rect 666 677 700 711
rect 666 609 700 643
rect 666 541 700 575
rect 666 473 700 507
rect 666 405 700 439
rect 666 337 700 371
rect 666 269 700 303
rect 666 201 700 235
<< psubdiff >>
rect 41 1187 111 1199
rect 41 1153 58 1187
rect 92 1153 111 1187
rect 41 1119 111 1153
rect 41 1085 58 1119
rect 92 1085 111 1119
rect 41 1051 111 1085
rect 41 1017 58 1051
rect 92 1017 111 1051
rect 41 983 111 1017
rect 41 949 58 983
rect 92 949 111 983
rect 41 915 111 949
rect 41 881 58 915
rect 92 881 111 915
rect 41 847 111 881
rect 41 813 58 847
rect 92 813 111 847
rect 41 779 111 813
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 715 1187 785 1199
rect 715 1153 734 1187
rect 768 1153 785 1187
rect 715 1119 785 1153
rect 715 1085 734 1119
rect 768 1085 785 1119
rect 715 1051 785 1085
rect 715 1017 734 1051
rect 768 1017 785 1051
rect 715 983 785 1017
rect 715 949 734 983
rect 768 949 785 983
rect 715 915 785 949
rect 715 881 734 915
rect 768 881 785 915
rect 715 847 785 881
rect 715 813 734 847
rect 768 813 785 847
rect 715 779 785 813
rect 715 745 734 779
rect 768 745 785 779
rect 715 711 785 745
rect 715 677 734 711
rect 768 677 785 711
rect 715 643 785 677
rect 715 609 734 643
rect 768 609 785 643
rect 715 575 785 609
rect 715 541 734 575
rect 768 541 785 575
rect 715 507 785 541
rect 715 473 734 507
rect 768 473 785 507
rect 715 439 785 473
rect 715 405 734 439
rect 768 405 785 439
rect 715 371 785 405
rect 715 337 734 371
rect 768 337 785 371
rect 715 303 785 337
rect 715 269 734 303
rect 768 269 785 303
rect 715 235 785 269
rect 715 201 734 235
rect 768 201 785 235
rect 715 189 785 201
<< psubdiffcont >>
rect 58 1153 92 1187
rect 58 1085 92 1119
rect 58 1017 92 1051
rect 58 949 92 983
rect 58 881 92 915
rect 58 813 92 847
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 734 1153 768 1187
rect 734 1085 768 1119
rect 734 1017 768 1051
rect 734 949 768 983
rect 734 881 768 915
rect 734 813 768 847
rect 734 745 768 779
rect 734 677 768 711
rect 734 609 768 643
rect 734 541 768 575
rect 734 473 768 507
rect 734 405 768 439
rect 734 337 768 371
rect 734 269 768 303
rect 734 201 768 235
<< poly >>
rect 243 1367 583 1388
rect 116 1275 201 1291
rect 116 1241 132 1275
rect 166 1241 201 1275
rect 243 1265 260 1367
rect 566 1265 583 1367
rect 243 1249 583 1265
rect 625 1275 710 1291
rect 116 1225 201 1241
rect 171 1199 201 1225
rect 257 1199 293 1249
rect 349 1199 385 1249
rect 441 1199 477 1249
rect 533 1199 569 1249
rect 625 1241 660 1275
rect 694 1241 710 1275
rect 625 1225 710 1241
rect 625 1199 655 1225
rect 171 163 201 189
rect 116 147 201 163
rect 116 113 132 147
rect 166 113 201 147
rect 257 139 293 189
rect 349 139 385 189
rect 441 139 477 189
rect 533 139 569 189
rect 625 163 655 189
rect 625 147 710 163
rect 116 97 201 113
rect 243 123 583 139
rect 243 21 260 123
rect 566 21 583 123
rect 625 113 660 147
rect 694 113 710 147
rect 625 97 710 113
rect 243 0 583 21
<< polycont >>
rect 132 1241 166 1275
rect 260 1265 566 1367
rect 660 1241 694 1275
rect 132 113 166 147
rect 260 21 566 123
rect 660 113 694 147
<< locali >>
rect 238 1369 588 1388
rect 116 1275 182 1291
rect 116 1241 132 1275
rect 166 1241 182 1275
rect 238 1263 252 1369
rect 574 1263 588 1369
rect 238 1249 588 1263
rect 644 1275 710 1291
rect 116 1225 182 1241
rect 644 1241 660 1275
rect 694 1241 710 1275
rect 644 1225 710 1241
rect 116 1203 160 1225
rect 666 1203 710 1225
rect 41 1187 160 1203
rect 41 1153 58 1187
rect 92 1179 126 1187
rect 94 1153 126 1179
rect 41 1145 60 1153
rect 94 1145 160 1153
rect 41 1119 160 1145
rect 41 1085 58 1119
rect 92 1107 126 1119
rect 94 1085 126 1107
rect 41 1073 60 1085
rect 94 1073 160 1085
rect 41 1051 160 1073
rect 41 1017 58 1051
rect 92 1035 126 1051
rect 94 1017 126 1035
rect 41 1001 60 1017
rect 94 1001 160 1017
rect 41 983 160 1001
rect 41 949 58 983
rect 92 963 126 983
rect 94 949 126 963
rect 41 929 60 949
rect 94 929 160 949
rect 41 915 160 929
rect 41 881 58 915
rect 92 891 126 915
rect 94 881 126 891
rect 41 857 60 881
rect 94 857 160 881
rect 41 847 160 857
rect 41 813 58 847
rect 92 819 126 847
rect 94 813 126 819
rect 41 785 60 813
rect 94 785 160 813
rect 41 779 160 785
rect 41 745 58 779
rect 92 747 126 779
rect 94 745 126 747
rect 41 713 60 745
rect 94 713 160 745
rect 41 711 160 713
rect 41 677 58 711
rect 92 677 126 711
rect 41 675 160 677
rect 41 643 60 675
rect 94 643 160 675
rect 41 609 58 643
rect 94 641 126 643
rect 92 609 126 641
rect 41 603 160 609
rect 41 575 60 603
rect 94 575 160 603
rect 41 541 58 575
rect 94 569 126 575
rect 92 541 126 569
rect 41 531 160 541
rect 41 507 60 531
rect 94 507 160 531
rect 41 473 58 507
rect 94 497 126 507
rect 92 473 126 497
rect 41 459 160 473
rect 41 439 60 459
rect 94 439 160 459
rect 41 405 58 439
rect 94 425 126 439
rect 92 405 126 425
rect 41 387 160 405
rect 41 371 60 387
rect 94 371 160 387
rect 41 337 58 371
rect 94 353 126 371
rect 92 337 126 353
rect 41 315 160 337
rect 41 303 60 315
rect 94 303 160 315
rect 41 269 58 303
rect 94 281 126 303
rect 92 269 126 281
rect 41 243 160 269
rect 41 235 60 243
rect 94 235 160 243
rect 41 201 58 235
rect 94 209 126 235
rect 92 201 126 209
rect 41 185 160 201
rect 212 1187 246 1203
rect 212 1119 246 1145
rect 212 1051 246 1073
rect 212 983 246 1001
rect 212 915 246 929
rect 212 847 246 857
rect 212 779 246 785
rect 212 711 246 713
rect 212 675 246 677
rect 212 603 246 609
rect 212 531 246 541
rect 212 459 246 473
rect 212 387 246 405
rect 212 315 246 337
rect 212 243 246 269
rect 212 185 246 201
rect 304 1187 338 1203
rect 304 1119 338 1145
rect 304 1051 338 1073
rect 304 983 338 1001
rect 304 915 338 929
rect 304 847 338 857
rect 304 779 338 785
rect 304 711 338 713
rect 304 675 338 677
rect 304 603 338 609
rect 304 531 338 541
rect 304 459 338 473
rect 304 387 338 405
rect 304 315 338 337
rect 304 243 338 269
rect 304 185 338 201
rect 396 1187 430 1203
rect 396 1119 430 1145
rect 396 1051 430 1073
rect 396 983 430 1001
rect 396 915 430 929
rect 396 847 430 857
rect 396 779 430 785
rect 396 711 430 713
rect 396 675 430 677
rect 396 603 430 609
rect 396 531 430 541
rect 396 459 430 473
rect 396 387 430 405
rect 396 315 430 337
rect 396 243 430 269
rect 396 185 430 201
rect 488 1187 522 1203
rect 488 1119 522 1145
rect 488 1051 522 1073
rect 488 983 522 1001
rect 488 915 522 929
rect 488 847 522 857
rect 488 779 522 785
rect 488 711 522 713
rect 488 675 522 677
rect 488 603 522 609
rect 488 531 522 541
rect 488 459 522 473
rect 488 387 522 405
rect 488 315 522 337
rect 488 243 522 269
rect 488 185 522 201
rect 580 1187 614 1203
rect 580 1119 614 1145
rect 580 1051 614 1073
rect 580 983 614 1001
rect 580 915 614 929
rect 580 847 614 857
rect 580 779 614 785
rect 580 711 614 713
rect 580 675 614 677
rect 580 603 614 609
rect 580 531 614 541
rect 580 459 614 473
rect 580 387 614 405
rect 580 315 614 337
rect 580 243 614 269
rect 580 185 614 201
rect 666 1187 785 1203
rect 700 1179 734 1187
rect 700 1153 732 1179
rect 768 1153 785 1187
rect 666 1145 732 1153
rect 766 1145 785 1153
rect 666 1119 785 1145
rect 700 1107 734 1119
rect 700 1085 732 1107
rect 768 1085 785 1119
rect 666 1073 732 1085
rect 766 1073 785 1085
rect 666 1051 785 1073
rect 700 1035 734 1051
rect 700 1017 732 1035
rect 768 1017 785 1051
rect 666 1001 732 1017
rect 766 1001 785 1017
rect 666 983 785 1001
rect 700 963 734 983
rect 700 949 732 963
rect 768 949 785 983
rect 666 929 732 949
rect 766 929 785 949
rect 666 915 785 929
rect 700 891 734 915
rect 700 881 732 891
rect 768 881 785 915
rect 666 857 732 881
rect 766 857 785 881
rect 666 847 785 857
rect 700 819 734 847
rect 700 813 732 819
rect 768 813 785 847
rect 666 785 732 813
rect 766 785 785 813
rect 666 779 785 785
rect 700 747 734 779
rect 700 745 732 747
rect 768 745 785 779
rect 666 713 732 745
rect 766 713 785 745
rect 666 711 785 713
rect 700 677 734 711
rect 768 677 785 711
rect 666 675 785 677
rect 666 643 732 675
rect 766 643 785 675
rect 700 641 732 643
rect 700 609 734 641
rect 768 609 785 643
rect 666 603 785 609
rect 666 575 732 603
rect 766 575 785 603
rect 700 569 732 575
rect 700 541 734 569
rect 768 541 785 575
rect 666 531 785 541
rect 666 507 732 531
rect 766 507 785 531
rect 700 497 732 507
rect 700 473 734 497
rect 768 473 785 507
rect 666 459 785 473
rect 666 439 732 459
rect 766 439 785 459
rect 700 425 732 439
rect 700 405 734 425
rect 768 405 785 439
rect 666 387 785 405
rect 666 371 732 387
rect 766 371 785 387
rect 700 353 732 371
rect 700 337 734 353
rect 768 337 785 371
rect 666 315 785 337
rect 666 303 732 315
rect 766 303 785 315
rect 700 281 732 303
rect 700 269 734 281
rect 768 269 785 303
rect 666 243 785 269
rect 666 235 732 243
rect 766 235 785 243
rect 700 209 732 235
rect 700 201 734 209
rect 768 201 785 235
rect 666 185 785 201
rect 116 163 160 185
rect 666 163 710 185
rect 116 147 182 163
rect 116 113 132 147
rect 166 113 182 147
rect 644 147 710 163
rect 116 97 182 113
rect 238 125 588 139
rect 238 19 252 125
rect 574 19 588 125
rect 644 113 660 147
rect 694 113 710 147
rect 644 97 710 113
rect 238 0 588 19
<< viali >>
rect 252 1367 574 1369
rect 252 1265 260 1367
rect 260 1265 566 1367
rect 566 1265 574 1367
rect 252 1263 574 1265
rect 60 1153 92 1179
rect 92 1153 94 1179
rect 60 1145 94 1153
rect 60 1085 92 1107
rect 92 1085 94 1107
rect 60 1073 94 1085
rect 60 1017 92 1035
rect 92 1017 94 1035
rect 60 1001 94 1017
rect 60 949 92 963
rect 92 949 94 963
rect 60 929 94 949
rect 60 881 92 891
rect 92 881 94 891
rect 60 857 94 881
rect 60 813 92 819
rect 92 813 94 819
rect 60 785 94 813
rect 60 745 92 747
rect 92 745 94 747
rect 60 713 94 745
rect 60 643 94 675
rect 60 641 92 643
rect 92 641 94 643
rect 60 575 94 603
rect 60 569 92 575
rect 92 569 94 575
rect 60 507 94 531
rect 60 497 92 507
rect 92 497 94 507
rect 60 439 94 459
rect 60 425 92 439
rect 92 425 94 439
rect 60 371 94 387
rect 60 353 92 371
rect 92 353 94 371
rect 60 303 94 315
rect 60 281 92 303
rect 92 281 94 303
rect 60 235 94 243
rect 60 209 92 235
rect 92 209 94 235
rect 212 1153 246 1179
rect 212 1145 246 1153
rect 212 1085 246 1107
rect 212 1073 246 1085
rect 212 1017 246 1035
rect 212 1001 246 1017
rect 212 949 246 963
rect 212 929 246 949
rect 212 881 246 891
rect 212 857 246 881
rect 212 813 246 819
rect 212 785 246 813
rect 212 745 246 747
rect 212 713 246 745
rect 212 643 246 675
rect 212 641 246 643
rect 212 575 246 603
rect 212 569 246 575
rect 212 507 246 531
rect 212 497 246 507
rect 212 439 246 459
rect 212 425 246 439
rect 212 371 246 387
rect 212 353 246 371
rect 212 303 246 315
rect 212 281 246 303
rect 212 235 246 243
rect 212 209 246 235
rect 304 1153 338 1179
rect 304 1145 338 1153
rect 304 1085 338 1107
rect 304 1073 338 1085
rect 304 1017 338 1035
rect 304 1001 338 1017
rect 304 949 338 963
rect 304 929 338 949
rect 304 881 338 891
rect 304 857 338 881
rect 304 813 338 819
rect 304 785 338 813
rect 304 745 338 747
rect 304 713 338 745
rect 304 643 338 675
rect 304 641 338 643
rect 304 575 338 603
rect 304 569 338 575
rect 304 507 338 531
rect 304 497 338 507
rect 304 439 338 459
rect 304 425 338 439
rect 304 371 338 387
rect 304 353 338 371
rect 304 303 338 315
rect 304 281 338 303
rect 304 235 338 243
rect 304 209 338 235
rect 396 1153 430 1179
rect 396 1145 430 1153
rect 396 1085 430 1107
rect 396 1073 430 1085
rect 396 1017 430 1035
rect 396 1001 430 1017
rect 396 949 430 963
rect 396 929 430 949
rect 396 881 430 891
rect 396 857 430 881
rect 396 813 430 819
rect 396 785 430 813
rect 396 745 430 747
rect 396 713 430 745
rect 396 643 430 675
rect 396 641 430 643
rect 396 575 430 603
rect 396 569 430 575
rect 396 507 430 531
rect 396 497 430 507
rect 396 439 430 459
rect 396 425 430 439
rect 396 371 430 387
rect 396 353 430 371
rect 396 303 430 315
rect 396 281 430 303
rect 396 235 430 243
rect 396 209 430 235
rect 488 1153 522 1179
rect 488 1145 522 1153
rect 488 1085 522 1107
rect 488 1073 522 1085
rect 488 1017 522 1035
rect 488 1001 522 1017
rect 488 949 522 963
rect 488 929 522 949
rect 488 881 522 891
rect 488 857 522 881
rect 488 813 522 819
rect 488 785 522 813
rect 488 745 522 747
rect 488 713 522 745
rect 488 643 522 675
rect 488 641 522 643
rect 488 575 522 603
rect 488 569 522 575
rect 488 507 522 531
rect 488 497 522 507
rect 488 439 522 459
rect 488 425 522 439
rect 488 371 522 387
rect 488 353 522 371
rect 488 303 522 315
rect 488 281 522 303
rect 488 235 522 243
rect 488 209 522 235
rect 580 1153 614 1179
rect 580 1145 614 1153
rect 580 1085 614 1107
rect 580 1073 614 1085
rect 580 1017 614 1035
rect 580 1001 614 1017
rect 580 949 614 963
rect 580 929 614 949
rect 580 881 614 891
rect 580 857 614 881
rect 580 813 614 819
rect 580 785 614 813
rect 580 745 614 747
rect 580 713 614 745
rect 580 643 614 675
rect 580 641 614 643
rect 580 575 614 603
rect 580 569 614 575
rect 580 507 614 531
rect 580 497 614 507
rect 580 439 614 459
rect 580 425 614 439
rect 580 371 614 387
rect 580 353 614 371
rect 580 303 614 315
rect 580 281 614 303
rect 580 235 614 243
rect 580 209 614 235
rect 732 1153 734 1179
rect 734 1153 766 1179
rect 732 1145 766 1153
rect 732 1085 734 1107
rect 734 1085 766 1107
rect 732 1073 766 1085
rect 732 1017 734 1035
rect 734 1017 766 1035
rect 732 1001 766 1017
rect 732 949 734 963
rect 734 949 766 963
rect 732 929 766 949
rect 732 881 734 891
rect 734 881 766 891
rect 732 857 766 881
rect 732 813 734 819
rect 734 813 766 819
rect 732 785 766 813
rect 732 745 734 747
rect 734 745 766 747
rect 732 713 766 745
rect 732 643 766 675
rect 732 641 734 643
rect 734 641 766 643
rect 732 575 766 603
rect 732 569 734 575
rect 734 569 766 575
rect 732 507 766 531
rect 732 497 734 507
rect 734 497 766 507
rect 732 439 766 459
rect 732 425 734 439
rect 734 425 766 439
rect 732 371 766 387
rect 732 353 734 371
rect 734 353 766 371
rect 732 303 766 315
rect 732 281 734 303
rect 734 281 766 303
rect 732 235 766 243
rect 732 209 734 235
rect 734 209 766 235
rect 252 123 574 125
rect 252 21 260 123
rect 260 21 566 123
rect 566 21 574 123
rect 252 19 574 21
<< metal1 >>
rect 236 1369 590 1388
rect 236 1263 252 1369
rect 574 1263 590 1369
rect 236 1251 590 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 203 1179 255 1191
rect 203 1145 212 1179
rect 246 1145 255 1179
rect 203 1107 255 1145
rect 203 1073 212 1107
rect 246 1073 255 1107
rect 203 1035 255 1073
rect 203 1001 212 1035
rect 246 1001 255 1035
rect 203 963 255 1001
rect 203 929 212 963
rect 246 929 255 963
rect 203 891 255 929
rect 203 857 212 891
rect 246 857 255 891
rect 203 819 255 857
rect 203 785 212 819
rect 246 785 255 819
rect 203 747 255 785
rect 203 713 212 747
rect 246 713 255 747
rect 203 675 255 713
rect 203 641 212 675
rect 246 641 255 675
rect 203 639 255 641
rect 203 575 212 587
rect 246 575 255 587
rect 203 511 212 523
rect 246 511 255 523
rect 203 447 212 459
rect 246 447 255 459
rect 203 387 255 395
rect 203 383 212 387
rect 246 383 255 387
rect 203 319 255 331
rect 203 255 255 267
rect 203 197 255 203
rect 295 1185 347 1191
rect 295 1121 347 1133
rect 295 1057 347 1069
rect 295 1001 304 1005
rect 338 1001 347 1005
rect 295 993 347 1001
rect 295 929 304 941
rect 338 929 347 941
rect 295 865 304 877
rect 338 865 347 877
rect 295 801 304 813
rect 338 801 347 813
rect 295 747 347 749
rect 295 713 304 747
rect 338 713 347 747
rect 295 675 347 713
rect 295 641 304 675
rect 338 641 347 675
rect 295 603 347 641
rect 295 569 304 603
rect 338 569 347 603
rect 295 531 347 569
rect 295 497 304 531
rect 338 497 347 531
rect 295 459 347 497
rect 295 425 304 459
rect 338 425 347 459
rect 295 387 347 425
rect 295 353 304 387
rect 338 353 347 387
rect 295 315 347 353
rect 295 281 304 315
rect 338 281 347 315
rect 295 243 347 281
rect 295 209 304 243
rect 338 209 347 243
rect 295 197 347 209
rect 387 1179 439 1191
rect 387 1145 396 1179
rect 430 1145 439 1179
rect 387 1107 439 1145
rect 387 1073 396 1107
rect 430 1073 439 1107
rect 387 1035 439 1073
rect 387 1001 396 1035
rect 430 1001 439 1035
rect 387 963 439 1001
rect 387 929 396 963
rect 430 929 439 963
rect 387 891 439 929
rect 387 857 396 891
rect 430 857 439 891
rect 387 819 439 857
rect 387 785 396 819
rect 430 785 439 819
rect 387 747 439 785
rect 387 713 396 747
rect 430 713 439 747
rect 387 675 439 713
rect 387 641 396 675
rect 430 641 439 675
rect 387 639 439 641
rect 387 575 396 587
rect 430 575 439 587
rect 387 511 396 523
rect 430 511 439 523
rect 387 447 396 459
rect 430 447 439 459
rect 387 387 439 395
rect 387 383 396 387
rect 430 383 439 387
rect 387 319 439 331
rect 387 255 439 267
rect 387 197 439 203
rect 479 1185 531 1191
rect 479 1121 531 1133
rect 479 1057 531 1069
rect 479 1001 488 1005
rect 522 1001 531 1005
rect 479 993 531 1001
rect 479 929 488 941
rect 522 929 531 941
rect 479 865 488 877
rect 522 865 531 877
rect 479 801 488 813
rect 522 801 531 813
rect 479 747 531 749
rect 479 713 488 747
rect 522 713 531 747
rect 479 675 531 713
rect 479 641 488 675
rect 522 641 531 675
rect 479 603 531 641
rect 479 569 488 603
rect 522 569 531 603
rect 479 531 531 569
rect 479 497 488 531
rect 522 497 531 531
rect 479 459 531 497
rect 479 425 488 459
rect 522 425 531 459
rect 479 387 531 425
rect 479 353 488 387
rect 522 353 531 387
rect 479 315 531 353
rect 479 281 488 315
rect 522 281 531 315
rect 479 243 531 281
rect 479 209 488 243
rect 522 209 531 243
rect 479 197 531 209
rect 571 1179 623 1191
rect 571 1145 580 1179
rect 614 1145 623 1179
rect 571 1107 623 1145
rect 571 1073 580 1107
rect 614 1073 623 1107
rect 571 1035 623 1073
rect 571 1001 580 1035
rect 614 1001 623 1035
rect 571 963 623 1001
rect 571 929 580 963
rect 614 929 623 963
rect 571 891 623 929
rect 571 857 580 891
rect 614 857 623 891
rect 571 819 623 857
rect 571 785 580 819
rect 614 785 623 819
rect 571 747 623 785
rect 571 713 580 747
rect 614 713 623 747
rect 571 675 623 713
rect 571 641 580 675
rect 614 641 623 675
rect 571 639 623 641
rect 571 575 580 587
rect 614 575 623 587
rect 571 511 580 523
rect 614 511 623 523
rect 571 447 580 459
rect 614 447 623 459
rect 571 387 623 395
rect 571 383 580 387
rect 614 383 623 387
rect 571 319 623 331
rect 571 255 623 267
rect 571 197 623 203
rect 726 1179 785 1191
rect 726 1145 732 1179
rect 766 1145 785 1179
rect 726 1107 785 1145
rect 726 1073 732 1107
rect 766 1073 785 1107
rect 726 1035 785 1073
rect 726 1001 732 1035
rect 766 1001 785 1035
rect 726 963 785 1001
rect 726 929 732 963
rect 766 929 785 963
rect 726 891 785 929
rect 726 857 732 891
rect 766 857 785 891
rect 726 819 785 857
rect 726 785 732 819
rect 766 785 785 819
rect 726 747 785 785
rect 726 713 732 747
rect 766 713 785 747
rect 726 675 785 713
rect 726 641 732 675
rect 766 641 785 675
rect 726 603 785 641
rect 726 569 732 603
rect 766 569 785 603
rect 726 531 785 569
rect 726 497 732 531
rect 766 497 785 531
rect 726 459 785 497
rect 726 425 732 459
rect 766 425 785 459
rect 726 387 785 425
rect 726 353 732 387
rect 766 353 785 387
rect 726 315 785 353
rect 726 281 732 315
rect 766 281 785 315
rect 726 243 785 281
rect 726 209 732 243
rect 766 209 785 243
rect 726 197 785 209
rect 236 125 590 137
rect 236 19 252 125
rect 574 19 590 125
rect 236 0 590 19
<< via1 >>
rect 203 603 255 639
rect 203 587 212 603
rect 212 587 246 603
rect 246 587 255 603
rect 203 569 212 575
rect 212 569 246 575
rect 246 569 255 575
rect 203 531 255 569
rect 203 523 212 531
rect 212 523 246 531
rect 246 523 255 531
rect 203 497 212 511
rect 212 497 246 511
rect 246 497 255 511
rect 203 459 255 497
rect 203 425 212 447
rect 212 425 246 447
rect 246 425 255 447
rect 203 395 255 425
rect 203 353 212 383
rect 212 353 246 383
rect 246 353 255 383
rect 203 331 255 353
rect 203 315 255 319
rect 203 281 212 315
rect 212 281 246 315
rect 246 281 255 315
rect 203 267 255 281
rect 203 243 255 255
rect 203 209 212 243
rect 212 209 246 243
rect 246 209 255 243
rect 203 203 255 209
rect 295 1179 347 1185
rect 295 1145 304 1179
rect 304 1145 338 1179
rect 338 1145 347 1179
rect 295 1133 347 1145
rect 295 1107 347 1121
rect 295 1073 304 1107
rect 304 1073 338 1107
rect 338 1073 347 1107
rect 295 1069 347 1073
rect 295 1035 347 1057
rect 295 1005 304 1035
rect 304 1005 338 1035
rect 338 1005 347 1035
rect 295 963 347 993
rect 295 941 304 963
rect 304 941 338 963
rect 338 941 347 963
rect 295 891 347 929
rect 295 877 304 891
rect 304 877 338 891
rect 338 877 347 891
rect 295 857 304 865
rect 304 857 338 865
rect 338 857 347 865
rect 295 819 347 857
rect 295 813 304 819
rect 304 813 338 819
rect 338 813 347 819
rect 295 785 304 801
rect 304 785 338 801
rect 338 785 347 801
rect 295 749 347 785
rect 387 603 439 639
rect 387 587 396 603
rect 396 587 430 603
rect 430 587 439 603
rect 387 569 396 575
rect 396 569 430 575
rect 430 569 439 575
rect 387 531 439 569
rect 387 523 396 531
rect 396 523 430 531
rect 430 523 439 531
rect 387 497 396 511
rect 396 497 430 511
rect 430 497 439 511
rect 387 459 439 497
rect 387 425 396 447
rect 396 425 430 447
rect 430 425 439 447
rect 387 395 439 425
rect 387 353 396 383
rect 396 353 430 383
rect 430 353 439 383
rect 387 331 439 353
rect 387 315 439 319
rect 387 281 396 315
rect 396 281 430 315
rect 430 281 439 315
rect 387 267 439 281
rect 387 243 439 255
rect 387 209 396 243
rect 396 209 430 243
rect 430 209 439 243
rect 387 203 439 209
rect 479 1179 531 1185
rect 479 1145 488 1179
rect 488 1145 522 1179
rect 522 1145 531 1179
rect 479 1133 531 1145
rect 479 1107 531 1121
rect 479 1073 488 1107
rect 488 1073 522 1107
rect 522 1073 531 1107
rect 479 1069 531 1073
rect 479 1035 531 1057
rect 479 1005 488 1035
rect 488 1005 522 1035
rect 522 1005 531 1035
rect 479 963 531 993
rect 479 941 488 963
rect 488 941 522 963
rect 522 941 531 963
rect 479 891 531 929
rect 479 877 488 891
rect 488 877 522 891
rect 522 877 531 891
rect 479 857 488 865
rect 488 857 522 865
rect 522 857 531 865
rect 479 819 531 857
rect 479 813 488 819
rect 488 813 522 819
rect 522 813 531 819
rect 479 785 488 801
rect 488 785 522 801
rect 522 785 531 801
rect 479 749 531 785
rect 571 603 623 639
rect 571 587 580 603
rect 580 587 614 603
rect 614 587 623 603
rect 571 569 580 575
rect 580 569 614 575
rect 614 569 623 575
rect 571 531 623 569
rect 571 523 580 531
rect 580 523 614 531
rect 614 523 623 531
rect 571 497 580 511
rect 580 497 614 511
rect 614 497 623 511
rect 571 459 623 497
rect 571 425 580 447
rect 580 425 614 447
rect 614 425 623 447
rect 571 395 623 425
rect 571 353 580 383
rect 580 353 614 383
rect 614 353 623 383
rect 571 331 623 353
rect 571 315 623 319
rect 571 281 580 315
rect 580 281 614 315
rect 614 281 623 315
rect 571 267 623 281
rect 571 243 623 255
rect 571 209 580 243
rect 580 209 614 243
rect 614 209 623 243
rect 571 203 623 209
<< metal2 >>
rect 14 1185 812 1191
rect 14 1133 295 1185
rect 347 1133 479 1185
rect 531 1133 812 1185
rect 14 1121 812 1133
rect 14 1069 295 1121
rect 347 1069 479 1121
rect 531 1069 812 1121
rect 14 1057 812 1069
rect 14 1005 295 1057
rect 347 1005 479 1057
rect 531 1005 812 1057
rect 14 993 812 1005
rect 14 941 295 993
rect 347 941 479 993
rect 531 941 812 993
rect 14 929 812 941
rect 14 877 295 929
rect 347 877 479 929
rect 531 877 812 929
rect 14 865 812 877
rect 14 813 295 865
rect 347 813 479 865
rect 531 813 812 865
rect 14 801 812 813
rect 14 749 295 801
rect 347 749 479 801
rect 531 749 812 801
rect 14 719 812 749
rect 14 639 812 669
rect 14 587 203 639
rect 255 587 387 639
rect 439 587 571 639
rect 623 587 812 639
rect 14 575 812 587
rect 14 523 203 575
rect 255 523 387 575
rect 439 523 571 575
rect 623 523 812 575
rect 14 511 812 523
rect 14 459 203 511
rect 255 459 387 511
rect 439 459 571 511
rect 623 459 812 511
rect 14 447 812 459
rect 14 395 203 447
rect 255 395 387 447
rect 439 395 571 447
rect 623 395 812 447
rect 14 383 812 395
rect 14 331 203 383
rect 255 331 387 383
rect 439 331 571 383
rect 623 331 812 383
rect 14 319 812 331
rect 14 267 203 319
rect 255 267 387 319
rect 439 267 571 319
rect 623 267 812 319
rect 14 255 812 267
rect 14 203 203 255
rect 255 203 387 255
rect 439 203 571 255
rect 623 203 812 255
rect 14 197 812 203
<< labels >>
flabel metal1 s 301 1286 535 1336 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 301 42 535 92 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 41 675 100 705 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 726 683 785 713 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel comment s 184 695 184 695 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 637 693 637 693 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 327 694 327 694 0 FreeSans 300 0 0 0 D
flabel comment s 241 694 241 694 0 FreeSans 300 0 0 0 S
flabel comment s 499 694 499 694 0 FreeSans 300 0 0 0 S
flabel comment s 413 694 413 694 0 FreeSans 300 0 0 0 S
flabel comment s 327 694 327 694 0 FreeSans 300 0 0 0 S
flabel comment s 241 694 241 694 0 FreeSans 300 0 0 0 S
flabel comment s 585 694 585 694 0 FreeSans 300 0 0 0 S
flabel comment s 499 694 499 694 0 FreeSans 300 0 0 0 D
flabel comment s 413 694 413 694 0 FreeSans 300 0 0 0 S
flabel metal2 s 14 384 35 512 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 908 35 1036 7 FreeSans 300 180 0 0 DRAIN
port 1 nsew
<< properties >>
string GDS_END 6431366
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6403244
string device primitive
<< end >>
