magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 1011 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 603 47 633 177
rect 687 47 717 177
rect 779 47 809 177
rect 864 47 894 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 603 297 633 497
rect 687 297 717 497
rect 779 297 809 497
rect 864 297 894 497
<< ndiff >>
rect 27 119 79 177
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 165 247 177
rect 193 131 203 165
rect 237 131 247 165
rect 193 47 247 131
rect 277 161 331 177
rect 277 127 287 161
rect 321 127 331 161
rect 277 93 331 127
rect 277 59 287 93
rect 321 59 331 93
rect 277 47 331 59
rect 361 109 415 177
rect 361 75 371 109
rect 405 75 415 109
rect 361 47 415 75
rect 445 93 497 177
rect 445 59 455 93
rect 489 59 497 93
rect 445 47 497 59
rect 551 93 603 177
rect 551 59 559 93
rect 593 59 603 93
rect 551 47 603 59
rect 633 165 687 177
rect 633 131 643 165
rect 677 131 687 165
rect 633 47 687 131
rect 717 93 779 177
rect 717 59 727 93
rect 761 59 779 93
rect 717 47 779 59
rect 809 165 864 177
rect 809 131 819 165
rect 853 131 864 165
rect 809 47 864 131
rect 894 93 985 177
rect 894 59 943 93
rect 977 59 985 93
rect 894 47 985 59
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 297 79 443
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 297 163 451
rect 193 401 247 497
rect 193 367 203 401
rect 237 367 247 401
rect 193 297 247 367
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 297 331 451
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 297 415 443
rect 445 485 497 497
rect 445 451 455 485
rect 489 451 497 485
rect 445 297 497 451
rect 551 485 603 497
rect 551 451 559 485
rect 593 451 603 485
rect 551 297 603 451
rect 633 343 687 497
rect 633 309 643 343
rect 677 309 687 343
rect 633 297 687 309
rect 717 485 779 497
rect 717 451 731 485
rect 765 451 779 485
rect 717 297 779 451
rect 809 417 864 497
rect 809 383 820 417
rect 854 383 864 417
rect 809 297 864 383
rect 894 485 985 497
rect 894 451 905 485
rect 939 451 985 485
rect 894 297 985 451
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 131 237 165
rect 287 127 321 161
rect 287 59 321 93
rect 371 75 405 109
rect 455 59 489 93
rect 559 59 593 93
rect 643 131 677 165
rect 727 59 761 93
rect 819 131 853 165
rect 943 59 977 93
<< pdiffc >>
rect 35 443 69 477
rect 119 451 153 485
rect 203 367 237 401
rect 287 451 321 485
rect 371 443 405 477
rect 455 451 489 485
rect 559 451 593 485
rect 643 309 677 343
rect 731 451 765 485
rect 820 383 854 417
rect 905 451 939 485
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 603 497 633 523
rect 687 497 717 523
rect 779 497 809 523
rect 864 497 894 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 415 265 445 297
rect 76 249 277 265
rect 76 215 86 249
rect 120 215 277 249
rect 76 199 277 215
rect 328 249 445 265
rect 603 265 633 297
rect 687 265 717 297
rect 779 265 809 297
rect 864 265 894 297
rect 603 259 724 265
rect 328 215 347 249
rect 381 215 445 249
rect 328 205 445 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 205
rect 415 177 445 205
rect 494 249 724 259
rect 494 215 510 249
rect 544 215 578 249
rect 612 215 646 249
rect 680 215 724 249
rect 494 199 724 215
rect 779 249 942 265
rect 779 215 893 249
rect 927 215 942 249
rect 779 199 942 215
rect 603 177 633 199
rect 687 177 717 199
rect 779 177 809 199
rect 864 177 894 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 603 21 633 47
rect 687 21 717 47
rect 779 21 809 47
rect 864 21 894 47
<< polycont >>
rect 86 215 120 249
rect 347 215 381 249
rect 510 215 544 249
rect 578 215 612 249
rect 646 215 680 249
rect 893 215 927 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 477 69 493
rect 17 443 35 477
rect 103 485 169 527
rect 103 451 119 485
rect 153 451 169 485
rect 271 485 337 527
rect 271 451 287 485
rect 321 451 337 485
rect 371 477 416 493
rect 17 427 69 443
rect 405 443 416 477
rect 371 427 416 443
rect 455 485 505 527
rect 489 451 505 485
rect 543 451 559 485
rect 593 451 731 485
rect 765 451 905 485
rect 939 451 995 485
rect 455 435 505 451
rect 17 333 52 427
rect 382 401 416 427
rect 543 401 820 417
rect 187 367 203 401
rect 237 367 347 401
rect 382 383 820 401
rect 854 383 870 417
rect 382 367 577 383
rect 313 333 347 367
rect 950 357 995 451
rect 627 333 643 343
rect 17 299 279 333
rect 313 309 643 333
rect 677 309 693 343
rect 313 299 693 309
rect 17 135 52 299
rect 245 265 279 299
rect 86 249 156 265
rect 120 215 156 249
rect 245 249 397 265
rect 245 231 347 249
rect 331 215 347 231
rect 381 215 397 249
rect 494 249 712 255
rect 494 215 510 249
rect 544 215 578 249
rect 612 215 646 249
rect 680 215 712 249
rect 862 249 927 323
rect 862 215 893 249
rect 86 199 156 215
rect 862 199 927 215
rect 116 145 156 199
rect 203 165 214 187
rect 248 153 251 187
rect 17 119 69 135
rect 17 85 35 119
rect 237 131 251 153
rect 203 115 251 131
rect 287 161 337 177
rect 321 127 337 161
rect 17 69 69 85
rect 103 93 167 109
rect 103 59 119 93
rect 153 59 167 93
rect 103 17 167 59
rect 287 93 337 127
rect 321 59 337 93
rect 371 165 693 181
rect 371 147 643 165
rect 371 109 405 147
rect 627 131 643 147
rect 677 131 693 165
rect 804 165 821 187
rect 804 153 819 165
rect 770 131 819 153
rect 853 131 869 165
rect 371 59 405 75
rect 455 93 489 109
rect 961 93 995 357
rect 543 59 559 93
rect 593 59 727 93
rect 761 59 943 93
rect 977 59 995 93
rect 287 17 337 59
rect 455 17 489 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 214 165 248 187
rect 214 153 237 165
rect 237 153 248 165
rect 770 153 804 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 202 187 260 193
rect 202 153 214 187
rect 248 184 260 187
rect 758 187 816 193
rect 758 184 770 187
rect 248 156 770 184
rect 248 153 260 156
rect 202 147 260 153
rect 758 153 770 156
rect 804 153 816 187
rect 758 147 816 153
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel locali s 950 425 984 459 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 862 289 896 323 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 862 221 896 255 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 950 357 984 391 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 494 221 528 255 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel locali s 586 221 620 255 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel locali s 678 221 712 255 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 mux2i_2
rlabel metal1 s 0 -48 1012 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_END 1705622
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1697608
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 25.300 0.000 
<< end >>
