magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__pfet_01v8__example_55959141808654  sky130_fd_pr__pfet_01v8__example_55959141808654_0
timestamp 1686671242
transform 0 -1 1756 1 0 197
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_55959141808654  sky130_fd_pr__pfet_01v8__example_55959141808654_1
timestamp 1686671242
transform 0 -1 3286 1 0 197
box -1 0 569 1
<< properties >>
string GDS_END 5685224
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 5653446
<< end >>
