magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< poly >>
rect 419 9430 579 9446
rect 419 9396 448 9430
rect 482 9396 516 9430
rect 550 9396 579 9430
rect -256 8806 -96 8822
rect -256 8772 -227 8806
rect -193 8772 -159 8806
rect -125 8772 -96 8806
rect 419 8162 448 8196
rect 482 8162 516 8196
rect 550 8162 579 8196
rect 419 8146 579 8162
rect 419 8088 579 8104
rect 419 8054 448 8088
rect 482 8054 516 8088
rect 550 8054 579 8088
rect 419 6820 448 6854
rect 482 6820 516 6854
rect 550 6820 579 6854
rect 419 6804 579 6820
rect -256 6338 -227 6372
rect -193 6338 -159 6372
rect -125 6338 -96 6372
rect -256 6322 -96 6338
rect -258 6080 -98 6096
rect -258 6046 -229 6080
rect -195 6046 -161 6080
rect -127 6046 -98 6080
rect -2 6080 158 6096
rect -2 6046 27 6080
rect 61 6046 95 6080
rect 129 6046 158 6080
<< polycont >>
rect 448 9396 482 9430
rect 516 9396 550 9430
rect -227 8772 -193 8806
rect -159 8772 -125 8806
rect 448 8162 482 8196
rect 516 8162 550 8196
rect 448 8054 482 8088
rect 516 8054 550 8088
rect 448 6820 482 6854
rect 516 6820 550 6854
rect -227 6338 -193 6372
rect -159 6338 -125 6372
rect -229 6046 -195 6080
rect -161 6046 -127 6080
rect 27 6046 61 6080
rect 95 6046 129 6080
<< npolyres >>
rect -256 6372 -96 8772
rect 419 8196 579 9396
rect 419 6854 579 8054
rect -258 1174 -98 6046
rect -2 1174 158 6046
rect -258 1014 158 1174
<< locali >>
rect 432 9396 448 9430
rect 482 9396 516 9430
rect 550 9396 566 9430
rect -243 8772 -227 8806
rect -193 8772 -159 8806
rect -125 8772 -109 8806
rect 432 8162 448 8196
rect 482 8162 516 8196
rect 550 8162 566 8196
rect 432 8054 448 8088
rect 482 8054 516 8088
rect 550 8054 566 8088
rect 432 6820 448 6854
rect 482 6820 516 6854
rect 550 6820 566 6854
rect -243 6338 -229 6372
rect -193 6338 -159 6372
rect -123 6338 -109 6372
rect -245 6046 -229 6080
rect -195 6046 -161 6080
rect -123 6046 -111 6080
rect 11 6046 27 6080
rect 61 6046 95 6080
rect 129 6046 145 6080
<< viali >>
rect -229 6338 -227 6372
rect -227 6338 -195 6372
rect -157 6338 -125 6372
rect -125 6338 -123 6372
rect -229 6046 -195 6080
rect -157 6046 -127 6080
rect -127 6046 -123 6080
<< metal1 >>
rect -241 6372 -111 6378
rect -241 6338 -229 6372
rect -195 6338 -157 6372
rect -123 6338 -111 6372
rect -241 6080 -111 6338
rect -241 6046 -229 6080
rect -195 6046 -157 6080
rect -123 6046 -111 6080
rect -241 6040 -111 6046
use sky130_fd_pr__res_bent_po__example_5595914180861  sky130_fd_pr__res_bent_po__example_5595914180861_0
timestamp 1686671242
transform 0 -1 -98 -1 0 6046
box -50 -243 -49 14
use sky130_fd_pr__res_bent_po__example_5595914180862  sky130_fd_pr__res_bent_po__example_5595914180862_0
timestamp 1686671242
transform 0 1 419 -1 0 9396
box -50 13 1185 14
use sky130_fd_pr__res_bent_po__example_5595914180862  sky130_fd_pr__res_bent_po__example_5595914180862_1
timestamp 1686671242
transform 0 1 419 -1 0 8054
box -50 13 1185 14
use sky130_fd_pr__res_bent_po__example_5595914180863  sky130_fd_pr__res_bent_po__example_5595914180863_0
timestamp 1686671242
transform 0 1 -256 -1 0 8772
box -50 13 2385 14
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1686671242
transform 1 0 -229 0 1 6338
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1686671242
transform 1 0 -229 0 1 6046
box 0 0 1 1
<< properties >>
string GDS_END 3731538
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3730974
<< end >>
