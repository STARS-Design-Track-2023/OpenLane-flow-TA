magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< locali >>
rect -4930 -2460 -4896 -2444
rect -4930 -2510 -4896 -2494
rect -4930 -3870 -4896 -3854
rect -4930 -3920 -4896 -3904
<< viali >>
rect -4930 -2494 -4896 -2460
rect -4930 -3904 -4896 -3870
<< metal1 >>
rect -4945 -2503 -4939 -2451
rect -4887 -2503 -4881 -2451
rect -4945 -3913 -4939 -3861
rect -4887 -3913 -4881 -3861
<< via1 >>
rect -4939 -2460 -4887 -2451
rect -4939 -2494 -4930 -2460
rect -4930 -2494 -4896 -2460
rect -4896 -2494 -4887 -2460
rect -4939 -2503 -4887 -2494
rect -4939 -3870 -4887 -3861
rect -4939 -3904 -4930 -3870
rect -4930 -3904 -4896 -3870
rect -4896 -3904 -4887 -3870
rect -4939 -3913 -4887 -3904
<< metal2 >>
rect -4941 -2449 -4885 -2440
rect -4941 -2514 -4885 -2505
rect -4526 -2449 -4470 -2440
rect -4526 -2514 -4470 -2505
rect -4512 -2679 -4484 -2514
rect -4526 -2688 -4470 -2679
rect -4526 -2753 -4470 -2744
rect -4662 -2812 -4606 -2803
rect -4662 -2877 -4606 -2868
rect -4648 -3850 -4620 -2877
rect -4941 -3859 -4885 -3850
rect -4941 -3924 -4885 -3915
rect -4662 -3859 -4606 -3850
rect -4662 -3924 -4606 -3915
<< via2 >>
rect -4941 -2451 -4885 -2449
rect -4941 -2503 -4939 -2451
rect -4939 -2503 -4887 -2451
rect -4887 -2503 -4885 -2451
rect -4941 -2505 -4885 -2503
rect -4526 -2505 -4470 -2449
rect -4526 -2744 -4470 -2688
rect -4662 -2868 -4606 -2812
rect -4941 -3861 -4885 -3859
rect -4941 -3913 -4939 -3861
rect -4939 -3913 -4887 -3861
rect -4887 -3913 -4885 -3861
rect -4941 -3915 -4885 -3913
rect -4662 -3915 -4606 -3859
<< metal3 >>
rect -4946 -2447 -4880 -2444
rect -4531 -2447 -4465 -2444
rect -4946 -2449 -4465 -2447
rect -4946 -2505 -4941 -2449
rect -4885 -2505 -4526 -2449
rect -4470 -2505 -4465 -2449
rect -4946 -2507 -4465 -2505
rect -4946 -2510 -4880 -2507
rect -4531 -2510 -4465 -2507
rect -4531 -2686 -4465 -2683
rect -4531 -2688 1278 -2686
rect -4531 -2744 -4526 -2688
rect -4470 -2744 1278 -2688
rect -4531 -2746 1278 -2744
rect -4531 -2749 -4465 -2746
rect -4667 -2810 -4601 -2807
rect -4667 -2812 1278 -2810
rect -4667 -2868 -4662 -2812
rect -4606 -2868 1278 -2812
rect -4667 -2870 1278 -2868
rect -4667 -2873 -4601 -2870
rect -4946 -3857 -4880 -3854
rect -4667 -3857 -4601 -3854
rect -4946 -3859 -4601 -3857
rect -4946 -3915 -4941 -3859
rect -4885 -3915 -4662 -3859
rect -4606 -3915 -4601 -3859
rect -4946 -3917 -4601 -3915
rect -4946 -3920 -4880 -3917
rect -4667 -3920 -4601 -3917
use contact_7  contact_7_0
timestamp 1686671242
transform 1 0 -4942 0 1 -2510
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1686671242
transform 1 0 -4942 0 1 -3920
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1686671242
transform 1 0 -4945 0 1 -2509
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1686671242
transform 1 0 -4945 0 1 -3919
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1686671242
transform 1 0 -4531 0 1 -2753
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1686671242
transform 1 0 -4946 0 1 -2514
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1686671242
transform 1 0 -4531 0 1 -2514
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1686671242
transform 1 0 -4667 0 1 -2877
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1686671242
transform 1 0 -4946 0 1 -3924
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1686671242
transform 1 0 -4667 0 1 -3924
box 0 0 1 1
<< properties >>
string FIXED_BBOX -4946 -3924 1278 -2440
string GDS_END 4888174
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4886934
<< end >>
