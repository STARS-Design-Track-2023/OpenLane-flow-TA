magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< metal4 >>
rect 0 34750 2000 39593
rect 0 13600 2000 18593
rect 0 12410 2000 13300
rect 0 11240 2000 12130
rect 0 10874 2000 10940
rect 0 10218 2000 10814
rect 0 9922 2000 10158
rect 0 9266 2000 9862
rect 0 9140 2000 9206
rect 0 7910 2000 8840
rect 0 6940 2000 7630
rect 0 5970 2000 6660
rect 0 4760 2000 5690
rect 0 3550 2000 4480
rect 0 2580 2000 3270
rect 0 1370 2000 2300
rect 0 0 2000 1090
<< metal5 >>
rect 0 34750 2000 39593
rect 0 13600 2000 18590
rect 0 12430 2000 13280
rect 0 11260 2000 12110
rect 0 9140 2000 10940
rect 0 7930 2000 8820
rect 0 6960 2000 7610
rect 0 5990 2000 6640
rect 0 4780 2000 5670
rect 0 3570 2000 4460
rect 0 2600 2000 3250
rect 0 1390 2000 2280
rect 0 20 2000 1070
<< labels >>
flabel metal4 s 1800 10218 2000 10814 0 FreeSans 800 0 0 0 AMUXBUS_A
port 1 nsew
flabel metal4 s 0 10218 200 10814 0 FreeSans 800 0 0 0 AMUXBUS_A
port 1 nsew
flabel metal4 s 1800 9266 2000 9862 0 FreeSans 800 0 0 0 AMUXBUS_B
port 2 nsew
flabel metal4 s 0 9266 200 9862 0 FreeSans 800 0 0 0 AMUXBUS_B
port 2 nsew
flabel metal4 s 1800 6940 2000 7630 0 FreeSans 800 0 0 0 VSSA
port 3 nsew
flabel metal5 s 1800 6960 2000 7610 0 FreeSans 800 0 0 0 VSSA
port 3 nsew
flabel metal4 s 1800 9140 2000 9206 0 FreeSans 800 0 0 0 VSSA
port 3 nsew
flabel metal4 s 1800 10874 2000 10940 0 FreeSans 800 0 0 0 VSSA
port 3 nsew
flabel metal5 s 1800 9140 2000 10940 0 FreeSans 800 0 0 0 VSSA
port 3 nsew
flabel metal4 s 0 6940 200 7630 0 FreeSans 800 0 0 0 VSSA
port 3 nsew
flabel metal5 s 0 6960 200 7610 0 FreeSans 800 0 0 0 VSSA
port 3 nsew
flabel metal4 s 0 9140 200 9206 0 FreeSans 800 0 0 0 VSSA
port 3 nsew
flabel metal4 s 0 10874 200 10940 0 FreeSans 800 0 0 0 VSSA
port 3 nsew
flabel metal5 s 0 9140 200 10940 0 FreeSans 800 0 0 0 VSSA
port 3 nsew
flabel metal4 s 1800 2580 2000 3270 0 FreeSans 800 0 0 0 VDDA
port 4 nsew
flabel metal5 s 1800 2600 2000 3250 0 FreeSans 800 0 0 0 VDDA
port 4 nsew
flabel metal4 s 0 2580 200 3270 0 FreeSans 800 0 0 0 VDDA
port 4 nsew
flabel metal5 s 0 2600 200 3250 0 FreeSans 800 0 0 0 VDDA
port 4 nsew
flabel metal4 s 1800 5970 2000 6660 0 FreeSans 800 0 0 0 VSWITCH
port 5 nsew
flabel metal5 s 1800 5990 2000 6640 0 FreeSans 800 0 0 0 VSWITCH
port 5 nsew
flabel metal4 s 0 5970 200 6660 0 FreeSans 800 0 0 0 VSWITCH
port 5 nsew
flabel metal5 s 0 5990 200 6640 0 FreeSans 800 0 0 0 VSWITCH
port 5 nsew
flabel metal4 s 1800 12410 2000 13300 0 FreeSans 800 0 0 0 VDDIO_Q
port 6 nsew
flabel metal5 s 1800 12430 2000 13280 0 FreeSans 800 0 0 0 VDDIO_Q
port 6 nsew
flabel metal4 s 0 12410 200 13300 0 FreeSans 800 0 0 0 VDDIO_Q
port 6 nsew
flabel metal5 s 0 12430 200 13280 0 FreeSans 800 0 0 0 VDDIO_Q
port 6 nsew
flabel metal4 s 1800 0 2000 1090 0 FreeSans 800 0 0 0 VCCHIB
port 7 nsew
flabel metal5 s 1800 20 2000 1070 0 FreeSans 800 0 0 0 VCCHIB
port 7 nsew
flabel metal4 s 0 0 200 1090 0 FreeSans 800 0 0 0 VCCHIB
port 7 nsew
flabel metal5 s 0 20 200 1070 0 FreeSans 800 0 0 0 VCCHIB
port 7 nsew
flabel metal4 s 1800 3550 2000 4480 0 FreeSans 800 0 0 0 VDDIO
port 8 nsew
flabel metal5 s 1800 3570 2000 4460 0 FreeSans 800 0 0 0 VDDIO
port 8 nsew
flabel metal4 s 1800 13600 2000 18593 0 FreeSans 800 0 0 0 VDDIO
port 8 nsew
flabel metal5 s 1800 13600 2000 18590 0 FreeSans 800 0 0 0 VDDIO
port 8 nsew
flabel metal4 s 0 3550 200 4480 0 FreeSans 800 0 0 0 VDDIO
port 8 nsew
flabel metal5 s 0 3570 200 4460 0 FreeSans 800 0 0 0 VDDIO
port 8 nsew
flabel metal4 s 0 13600 200 18593 0 FreeSans 800 0 0 0 VDDIO
port 8 nsew
flabel metal5 s 0 13600 200 18590 0 FreeSans 800 0 0 0 VDDIO
port 8 nsew
flabel metal4 s 1800 1370 2000 2300 0 FreeSans 800 0 0 0 VCCD
port 9 nsew
flabel metal5 s 1800 1390 2000 2280 0 FreeSans 800 0 0 0 VCCD
port 9 nsew
flabel metal4 s 0 1370 200 2300 0 FreeSans 800 0 0 0 VCCD
port 9 nsew
flabel metal5 s 0 1390 200 2280 0 FreeSans 800 0 0 0 VCCD
port 9 nsew
flabel metal5 s 1800 34750 2000 39593 0 FreeSans 800 0 0 0 VSSIO
port 10 nsew
flabel metal4 s 1800 4760 2000 5690 0 FreeSans 800 0 0 0 VSSIO
port 10 nsew
flabel metal5 s 1800 4780 2000 5670 0 FreeSans 800 0 0 0 VSSIO
port 10 nsew
flabel metal5 s 0 34750 200 39593 0 FreeSans 800 0 0 0 VSSIO
port 10 nsew
flabel metal4 s 0 4760 200 5690 0 FreeSans 800 0 0 0 VSSIO
port 10 nsew
flabel metal5 s 0 4780 200 5670 0 FreeSans 800 0 0 0 VSSIO
port 10 nsew
flabel metal4 s 1800 7910 2000 8840 0 FreeSans 800 0 0 0 VSSD
port 11 nsew
flabel metal5 s 1800 7930 2000 8820 0 FreeSans 800 0 0 0 VSSD
port 11 nsew
flabel metal4 s 0 7910 200 8840 0 FreeSans 800 0 0 0 VSSD
port 11 nsew
flabel metal5 s 0 7930 200 8820 0 FreeSans 800 0 0 0 VSSD
port 11 nsew
flabel metal4 s 1800 11240 2000 12130 0 FreeSans 800 0 0 0 VSSIO_Q
port 12 nsew
flabel metal5 s 1800 11260 2000 12110 0 FreeSans 800 0 0 0 VSSIO_Q
port 12 nsew
flabel metal4 s 0 11240 200 12130 0 FreeSans 800 0 0 0 VSSIO_Q
port 12 nsew
flabel metal5 s 0 11260 200 12110 0 FreeSans 800 0 0 0 VSSIO_Q
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 2000 39593
string GDS_END 3752122
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 3742858
<< end >>
