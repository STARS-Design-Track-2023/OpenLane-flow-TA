magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< poly >>
rect 0 2322 11146 2338
rect 0 2288 34 2322
rect 68 2288 102 2322
rect 136 2288 170 2322
rect 204 2288 238 2322
rect 272 2288 306 2322
rect 340 2288 374 2322
rect 408 2288 442 2322
rect 476 2288 510 2322
rect 544 2288 578 2322
rect 612 2288 646 2322
rect 680 2288 714 2322
rect 748 2288 782 2322
rect 816 2288 850 2322
rect 884 2288 918 2322
rect 952 2288 986 2322
rect 1020 2288 1054 2322
rect 1088 2288 1122 2322
rect 1156 2288 1190 2322
rect 1224 2288 1258 2322
rect 1292 2288 1326 2322
rect 1360 2288 1394 2322
rect 1428 2288 1462 2322
rect 1496 2288 1530 2322
rect 1564 2288 1598 2322
rect 1632 2288 1666 2322
rect 1700 2288 1734 2322
rect 1768 2288 1802 2322
rect 1836 2288 1870 2322
rect 1904 2288 1938 2322
rect 1972 2288 2006 2322
rect 2040 2288 2074 2322
rect 2108 2288 2142 2322
rect 2176 2288 2210 2322
rect 2244 2288 2278 2322
rect 2312 2288 2346 2322
rect 2380 2288 2414 2322
rect 2448 2288 2482 2322
rect 2516 2288 2550 2322
rect 2584 2288 2618 2322
rect 2652 2288 2686 2322
rect 2720 2288 2754 2322
rect 2788 2288 2822 2322
rect 2856 2288 2890 2322
rect 2924 2288 2958 2322
rect 2992 2288 3026 2322
rect 3060 2288 3094 2322
rect 3128 2288 3162 2322
rect 3196 2288 3230 2322
rect 3264 2288 3298 2322
rect 3332 2288 3366 2322
rect 3400 2288 3434 2322
rect 3468 2288 3502 2322
rect 3536 2288 3570 2322
rect 3604 2288 3638 2322
rect 3672 2288 3706 2322
rect 3740 2288 3774 2322
rect 3808 2288 3842 2322
rect 3876 2288 3910 2322
rect 3944 2288 3978 2322
rect 4012 2288 4046 2322
rect 4080 2288 4114 2322
rect 4148 2288 4182 2322
rect 4216 2288 4250 2322
rect 4284 2288 4318 2322
rect 4352 2288 4386 2322
rect 4420 2288 4454 2322
rect 4488 2288 4522 2322
rect 4556 2288 4590 2322
rect 4624 2288 4658 2322
rect 4692 2288 4726 2322
rect 4760 2288 4794 2322
rect 4828 2288 4862 2322
rect 4896 2288 4930 2322
rect 4964 2288 4998 2322
rect 5032 2288 5066 2322
rect 5100 2288 5134 2322
rect 5168 2288 5202 2322
rect 5236 2288 5270 2322
rect 5304 2288 5338 2322
rect 5372 2288 5406 2322
rect 5440 2288 5474 2322
rect 5508 2288 5542 2322
rect 5576 2288 5610 2322
rect 5644 2288 5678 2322
rect 5712 2288 5746 2322
rect 5780 2288 5814 2322
rect 5848 2288 5882 2322
rect 5916 2288 5950 2322
rect 5984 2288 6018 2322
rect 6052 2288 6086 2322
rect 6120 2288 6154 2322
rect 6188 2288 6222 2322
rect 6256 2288 6290 2322
rect 6324 2288 6358 2322
rect 6392 2288 6426 2322
rect 6460 2288 6494 2322
rect 6528 2288 6562 2322
rect 6596 2288 6630 2322
rect 6664 2288 6698 2322
rect 6732 2288 6766 2322
rect 6800 2288 6834 2322
rect 6868 2288 6902 2322
rect 6936 2288 6970 2322
rect 7004 2288 7038 2322
rect 7072 2288 7106 2322
rect 7140 2288 7174 2322
rect 7208 2288 7242 2322
rect 7276 2288 7310 2322
rect 7344 2288 7378 2322
rect 7412 2288 7446 2322
rect 7480 2288 7514 2322
rect 7548 2288 7582 2322
rect 7616 2288 7650 2322
rect 7684 2288 7718 2322
rect 7752 2288 7786 2322
rect 7820 2288 7854 2322
rect 7888 2288 7922 2322
rect 7956 2288 7990 2322
rect 8024 2288 8058 2322
rect 8092 2288 8126 2322
rect 8160 2288 8194 2322
rect 8228 2288 8262 2322
rect 8296 2288 8330 2322
rect 8364 2288 8398 2322
rect 8432 2288 8466 2322
rect 8500 2288 8534 2322
rect 8568 2288 8602 2322
rect 8636 2288 8670 2322
rect 8704 2288 8738 2322
rect 8772 2288 8806 2322
rect 8840 2288 8874 2322
rect 8908 2288 8942 2322
rect 8976 2288 9010 2322
rect 9044 2288 9078 2322
rect 9112 2288 9146 2322
rect 9180 2288 9214 2322
rect 9248 2288 9282 2322
rect 9316 2288 9350 2322
rect 9384 2288 9418 2322
rect 9452 2288 9486 2322
rect 9520 2288 9554 2322
rect 9588 2288 9622 2322
rect 9656 2288 9690 2322
rect 9724 2288 9758 2322
rect 9792 2288 9826 2322
rect 9860 2288 9894 2322
rect 9928 2288 9962 2322
rect 9996 2288 10030 2322
rect 10064 2288 10098 2322
rect 10132 2288 10166 2322
rect 10200 2288 10234 2322
rect 10268 2288 10302 2322
rect 10336 2288 10370 2322
rect 10404 2288 10438 2322
rect 10472 2288 10506 2322
rect 10540 2288 10574 2322
rect 10608 2288 10642 2322
rect 10676 2288 10710 2322
rect 10744 2288 10778 2322
rect 10812 2288 10846 2322
rect 10880 2288 10914 2322
rect 10948 2288 10982 2322
rect 11016 2288 11050 2322
rect 11084 2288 11146 2322
rect 0 2272 11146 2288
rect 0 108 30 2272
rect 72 66 102 2230
rect 144 108 174 2272
rect 216 66 246 2230
rect 288 108 318 2272
rect 360 66 390 2230
rect 432 108 462 2272
rect 504 66 534 2230
rect 576 108 606 2272
rect 648 66 678 2230
rect 720 108 750 2272
rect 792 66 822 2230
rect 864 108 894 2272
rect 936 66 966 2230
rect 1008 108 1038 2272
rect 1080 66 1110 2230
rect 1152 108 1182 2272
rect 1224 66 1254 2230
rect 1296 108 1326 2272
rect 1368 66 1398 2230
rect 1440 108 1470 2272
rect 1512 66 1542 2230
rect 1584 108 1614 2272
rect 1656 66 1686 2230
rect 1728 108 1758 2272
rect 1800 66 1830 2230
rect 1872 108 1902 2272
rect 1944 66 1974 2230
rect 2016 108 2046 2272
rect 2088 66 2118 2230
rect 2160 108 2190 2272
rect 2232 66 2262 2230
rect 2304 108 2334 2272
rect 2376 66 2406 2230
rect 2448 108 2478 2272
rect 2520 66 2550 2230
rect 2592 108 2622 2272
rect 2664 66 2694 2230
rect 2736 108 2766 2272
rect 2808 66 2838 2230
rect 2880 108 2910 2272
rect 2952 66 2982 2230
rect 3024 108 3054 2272
rect 3096 66 3126 2230
rect 3168 108 3198 2272
rect 3240 66 3270 2230
rect 3312 108 3342 2272
rect 3384 66 3414 2230
rect 3456 108 3486 2272
rect 3528 66 3558 2230
rect 3600 108 3630 2272
rect 3672 66 3702 2230
rect 3744 108 3774 2272
rect 3816 66 3846 2230
rect 3888 108 3918 2272
rect 3960 66 3990 2230
rect 4032 108 4062 2272
rect 4104 66 4134 2230
rect 4176 108 4206 2272
rect 4248 66 4278 2230
rect 4320 108 4350 2272
rect 4392 66 4422 2230
rect 4464 108 4494 2272
rect 4536 66 4566 2230
rect 4608 108 4638 2272
rect 4680 66 4710 2230
rect 4752 108 4782 2272
rect 4824 66 4854 2230
rect 4896 108 4926 2272
rect 4968 66 4998 2230
rect 5040 108 5070 2272
rect 5112 66 5142 2230
rect 5184 108 5214 2272
rect 5256 66 5286 2230
rect 5328 108 5358 2272
rect 5400 66 5430 2230
rect 5472 108 5502 2272
rect 5544 66 5574 2230
rect 5616 108 5646 2272
rect 5688 66 5718 2230
rect 5760 108 5790 2272
rect 5832 66 5862 2230
rect 5904 108 5934 2272
rect 5976 66 6006 2230
rect 6048 108 6078 2272
rect 6120 66 6150 2230
rect 6192 108 6222 2272
rect 6264 66 6294 2230
rect 6336 108 6366 2272
rect 6408 66 6438 2230
rect 6480 108 6510 2272
rect 6552 66 6582 2230
rect 6624 108 6654 2272
rect 6696 66 6726 2230
rect 6768 108 6798 2272
rect 6840 66 6870 2230
rect 6912 108 6942 2272
rect 6984 66 7014 2230
rect 7056 108 7086 2272
rect 7128 66 7158 2230
rect 7200 108 7230 2272
rect 7272 66 7302 2230
rect 7344 108 7374 2272
rect 7416 66 7446 2230
rect 7488 108 7518 2272
rect 7560 66 7590 2230
rect 7632 108 7662 2272
rect 7704 66 7734 2230
rect 7776 108 7806 2272
rect 7848 66 7878 2230
rect 7920 108 7950 2272
rect 7992 66 8022 2230
rect 8064 108 8094 2272
rect 8136 66 8166 2230
rect 8208 108 8238 2272
rect 8280 66 8310 2230
rect 8352 108 8382 2272
rect 8424 66 8454 2230
rect 8496 108 8526 2272
rect 8568 66 8598 2230
rect 8640 108 8670 2272
rect 8712 66 8742 2230
rect 8784 108 8814 2272
rect 8856 66 8886 2230
rect 8928 108 8958 2272
rect 9000 66 9030 2230
rect 9072 108 9102 2272
rect 9144 66 9174 2230
rect 9216 108 9246 2272
rect 9288 66 9318 2230
rect 9360 108 9390 2272
rect 9432 66 9462 2230
rect 9504 108 9534 2272
rect 9576 66 9606 2230
rect 9648 108 9678 2272
rect 9720 66 9750 2230
rect 9792 108 9822 2272
rect 9864 66 9894 2230
rect 9936 108 9966 2272
rect 10008 66 10038 2230
rect 10080 108 10110 2272
rect 10152 66 10182 2230
rect 10224 108 10254 2272
rect 10296 66 10326 2230
rect 10368 108 10398 2272
rect 10440 66 10470 2230
rect 10512 108 10542 2272
rect 10584 66 10614 2230
rect 10656 108 10686 2272
rect 10728 66 10758 2230
rect 10800 108 10830 2272
rect 10872 66 10902 2230
rect 10944 108 10974 2272
rect 11016 66 11046 2230
rect 11088 108 11146 2272
rect 0 50 11146 66
rect 0 16 34 50
rect 68 16 102 50
rect 136 16 170 50
rect 204 16 238 50
rect 272 16 306 50
rect 340 16 374 50
rect 408 16 442 50
rect 476 16 510 50
rect 544 16 578 50
rect 612 16 646 50
rect 680 16 714 50
rect 748 16 782 50
rect 816 16 850 50
rect 884 16 918 50
rect 952 16 986 50
rect 1020 16 1054 50
rect 1088 16 1122 50
rect 1156 16 1190 50
rect 1224 16 1258 50
rect 1292 16 1326 50
rect 1360 16 1394 50
rect 1428 16 1462 50
rect 1496 16 1530 50
rect 1564 16 1598 50
rect 1632 16 1666 50
rect 1700 16 1734 50
rect 1768 16 1802 50
rect 1836 16 1870 50
rect 1904 16 1938 50
rect 1972 16 2006 50
rect 2040 16 2074 50
rect 2108 16 2142 50
rect 2176 16 2210 50
rect 2244 16 2278 50
rect 2312 16 2346 50
rect 2380 16 2414 50
rect 2448 16 2482 50
rect 2516 16 2550 50
rect 2584 16 2618 50
rect 2652 16 2686 50
rect 2720 16 2754 50
rect 2788 16 2822 50
rect 2856 16 2890 50
rect 2924 16 2958 50
rect 2992 16 3026 50
rect 3060 16 3094 50
rect 3128 16 3162 50
rect 3196 16 3230 50
rect 3264 16 3298 50
rect 3332 16 3366 50
rect 3400 16 3434 50
rect 3468 16 3502 50
rect 3536 16 3570 50
rect 3604 16 3638 50
rect 3672 16 3706 50
rect 3740 16 3774 50
rect 3808 16 3842 50
rect 3876 16 3910 50
rect 3944 16 3978 50
rect 4012 16 4046 50
rect 4080 16 4114 50
rect 4148 16 4182 50
rect 4216 16 4250 50
rect 4284 16 4318 50
rect 4352 16 4386 50
rect 4420 16 4454 50
rect 4488 16 4522 50
rect 4556 16 4590 50
rect 4624 16 4658 50
rect 4692 16 4726 50
rect 4760 16 4794 50
rect 4828 16 4862 50
rect 4896 16 4930 50
rect 4964 16 4998 50
rect 5032 16 5066 50
rect 5100 16 5134 50
rect 5168 16 5202 50
rect 5236 16 5270 50
rect 5304 16 5338 50
rect 5372 16 5406 50
rect 5440 16 5474 50
rect 5508 16 5542 50
rect 5576 16 5610 50
rect 5644 16 5678 50
rect 5712 16 5746 50
rect 5780 16 5814 50
rect 5848 16 5882 50
rect 5916 16 5950 50
rect 5984 16 6018 50
rect 6052 16 6086 50
rect 6120 16 6154 50
rect 6188 16 6222 50
rect 6256 16 6290 50
rect 6324 16 6358 50
rect 6392 16 6426 50
rect 6460 16 6494 50
rect 6528 16 6562 50
rect 6596 16 6630 50
rect 6664 16 6698 50
rect 6732 16 6766 50
rect 6800 16 6834 50
rect 6868 16 6902 50
rect 6936 16 6970 50
rect 7004 16 7038 50
rect 7072 16 7106 50
rect 7140 16 7174 50
rect 7208 16 7242 50
rect 7276 16 7310 50
rect 7344 16 7378 50
rect 7412 16 7446 50
rect 7480 16 7514 50
rect 7548 16 7582 50
rect 7616 16 7650 50
rect 7684 16 7718 50
rect 7752 16 7786 50
rect 7820 16 7854 50
rect 7888 16 7922 50
rect 7956 16 7990 50
rect 8024 16 8058 50
rect 8092 16 8126 50
rect 8160 16 8194 50
rect 8228 16 8262 50
rect 8296 16 8330 50
rect 8364 16 8398 50
rect 8432 16 8466 50
rect 8500 16 8534 50
rect 8568 16 8602 50
rect 8636 16 8670 50
rect 8704 16 8738 50
rect 8772 16 8806 50
rect 8840 16 8874 50
rect 8908 16 8942 50
rect 8976 16 9010 50
rect 9044 16 9078 50
rect 9112 16 9146 50
rect 9180 16 9214 50
rect 9248 16 9282 50
rect 9316 16 9350 50
rect 9384 16 9418 50
rect 9452 16 9486 50
rect 9520 16 9554 50
rect 9588 16 9622 50
rect 9656 16 9690 50
rect 9724 16 9758 50
rect 9792 16 9826 50
rect 9860 16 9894 50
rect 9928 16 9962 50
rect 9996 16 10030 50
rect 10064 16 10098 50
rect 10132 16 10166 50
rect 10200 16 10234 50
rect 10268 16 10302 50
rect 10336 16 10370 50
rect 10404 16 10438 50
rect 10472 16 10506 50
rect 10540 16 10574 50
rect 10608 16 10642 50
rect 10676 16 10710 50
rect 10744 16 10778 50
rect 10812 16 10846 50
rect 10880 16 10914 50
rect 10948 16 10982 50
rect 11016 16 11050 50
rect 11084 16 11146 50
rect 0 0 11146 16
<< polycont >>
rect 34 2288 68 2322
rect 102 2288 136 2322
rect 170 2288 204 2322
rect 238 2288 272 2322
rect 306 2288 340 2322
rect 374 2288 408 2322
rect 442 2288 476 2322
rect 510 2288 544 2322
rect 578 2288 612 2322
rect 646 2288 680 2322
rect 714 2288 748 2322
rect 782 2288 816 2322
rect 850 2288 884 2322
rect 918 2288 952 2322
rect 986 2288 1020 2322
rect 1054 2288 1088 2322
rect 1122 2288 1156 2322
rect 1190 2288 1224 2322
rect 1258 2288 1292 2322
rect 1326 2288 1360 2322
rect 1394 2288 1428 2322
rect 1462 2288 1496 2322
rect 1530 2288 1564 2322
rect 1598 2288 1632 2322
rect 1666 2288 1700 2322
rect 1734 2288 1768 2322
rect 1802 2288 1836 2322
rect 1870 2288 1904 2322
rect 1938 2288 1972 2322
rect 2006 2288 2040 2322
rect 2074 2288 2108 2322
rect 2142 2288 2176 2322
rect 2210 2288 2244 2322
rect 2278 2288 2312 2322
rect 2346 2288 2380 2322
rect 2414 2288 2448 2322
rect 2482 2288 2516 2322
rect 2550 2288 2584 2322
rect 2618 2288 2652 2322
rect 2686 2288 2720 2322
rect 2754 2288 2788 2322
rect 2822 2288 2856 2322
rect 2890 2288 2924 2322
rect 2958 2288 2992 2322
rect 3026 2288 3060 2322
rect 3094 2288 3128 2322
rect 3162 2288 3196 2322
rect 3230 2288 3264 2322
rect 3298 2288 3332 2322
rect 3366 2288 3400 2322
rect 3434 2288 3468 2322
rect 3502 2288 3536 2322
rect 3570 2288 3604 2322
rect 3638 2288 3672 2322
rect 3706 2288 3740 2322
rect 3774 2288 3808 2322
rect 3842 2288 3876 2322
rect 3910 2288 3944 2322
rect 3978 2288 4012 2322
rect 4046 2288 4080 2322
rect 4114 2288 4148 2322
rect 4182 2288 4216 2322
rect 4250 2288 4284 2322
rect 4318 2288 4352 2322
rect 4386 2288 4420 2322
rect 4454 2288 4488 2322
rect 4522 2288 4556 2322
rect 4590 2288 4624 2322
rect 4658 2288 4692 2322
rect 4726 2288 4760 2322
rect 4794 2288 4828 2322
rect 4862 2288 4896 2322
rect 4930 2288 4964 2322
rect 4998 2288 5032 2322
rect 5066 2288 5100 2322
rect 5134 2288 5168 2322
rect 5202 2288 5236 2322
rect 5270 2288 5304 2322
rect 5338 2288 5372 2322
rect 5406 2288 5440 2322
rect 5474 2288 5508 2322
rect 5542 2288 5576 2322
rect 5610 2288 5644 2322
rect 5678 2288 5712 2322
rect 5746 2288 5780 2322
rect 5814 2288 5848 2322
rect 5882 2288 5916 2322
rect 5950 2288 5984 2322
rect 6018 2288 6052 2322
rect 6086 2288 6120 2322
rect 6154 2288 6188 2322
rect 6222 2288 6256 2322
rect 6290 2288 6324 2322
rect 6358 2288 6392 2322
rect 6426 2288 6460 2322
rect 6494 2288 6528 2322
rect 6562 2288 6596 2322
rect 6630 2288 6664 2322
rect 6698 2288 6732 2322
rect 6766 2288 6800 2322
rect 6834 2288 6868 2322
rect 6902 2288 6936 2322
rect 6970 2288 7004 2322
rect 7038 2288 7072 2322
rect 7106 2288 7140 2322
rect 7174 2288 7208 2322
rect 7242 2288 7276 2322
rect 7310 2288 7344 2322
rect 7378 2288 7412 2322
rect 7446 2288 7480 2322
rect 7514 2288 7548 2322
rect 7582 2288 7616 2322
rect 7650 2288 7684 2322
rect 7718 2288 7752 2322
rect 7786 2288 7820 2322
rect 7854 2288 7888 2322
rect 7922 2288 7956 2322
rect 7990 2288 8024 2322
rect 8058 2288 8092 2322
rect 8126 2288 8160 2322
rect 8194 2288 8228 2322
rect 8262 2288 8296 2322
rect 8330 2288 8364 2322
rect 8398 2288 8432 2322
rect 8466 2288 8500 2322
rect 8534 2288 8568 2322
rect 8602 2288 8636 2322
rect 8670 2288 8704 2322
rect 8738 2288 8772 2322
rect 8806 2288 8840 2322
rect 8874 2288 8908 2322
rect 8942 2288 8976 2322
rect 9010 2288 9044 2322
rect 9078 2288 9112 2322
rect 9146 2288 9180 2322
rect 9214 2288 9248 2322
rect 9282 2288 9316 2322
rect 9350 2288 9384 2322
rect 9418 2288 9452 2322
rect 9486 2288 9520 2322
rect 9554 2288 9588 2322
rect 9622 2288 9656 2322
rect 9690 2288 9724 2322
rect 9758 2288 9792 2322
rect 9826 2288 9860 2322
rect 9894 2288 9928 2322
rect 9962 2288 9996 2322
rect 10030 2288 10064 2322
rect 10098 2288 10132 2322
rect 10166 2288 10200 2322
rect 10234 2288 10268 2322
rect 10302 2288 10336 2322
rect 10370 2288 10404 2322
rect 10438 2288 10472 2322
rect 10506 2288 10540 2322
rect 10574 2288 10608 2322
rect 10642 2288 10676 2322
rect 10710 2288 10744 2322
rect 10778 2288 10812 2322
rect 10846 2288 10880 2322
rect 10914 2288 10948 2322
rect 10982 2288 11016 2322
rect 11050 2288 11084 2322
rect 34 16 68 50
rect 102 16 136 50
rect 170 16 204 50
rect 238 16 272 50
rect 306 16 340 50
rect 374 16 408 50
rect 442 16 476 50
rect 510 16 544 50
rect 578 16 612 50
rect 646 16 680 50
rect 714 16 748 50
rect 782 16 816 50
rect 850 16 884 50
rect 918 16 952 50
rect 986 16 1020 50
rect 1054 16 1088 50
rect 1122 16 1156 50
rect 1190 16 1224 50
rect 1258 16 1292 50
rect 1326 16 1360 50
rect 1394 16 1428 50
rect 1462 16 1496 50
rect 1530 16 1564 50
rect 1598 16 1632 50
rect 1666 16 1700 50
rect 1734 16 1768 50
rect 1802 16 1836 50
rect 1870 16 1904 50
rect 1938 16 1972 50
rect 2006 16 2040 50
rect 2074 16 2108 50
rect 2142 16 2176 50
rect 2210 16 2244 50
rect 2278 16 2312 50
rect 2346 16 2380 50
rect 2414 16 2448 50
rect 2482 16 2516 50
rect 2550 16 2584 50
rect 2618 16 2652 50
rect 2686 16 2720 50
rect 2754 16 2788 50
rect 2822 16 2856 50
rect 2890 16 2924 50
rect 2958 16 2992 50
rect 3026 16 3060 50
rect 3094 16 3128 50
rect 3162 16 3196 50
rect 3230 16 3264 50
rect 3298 16 3332 50
rect 3366 16 3400 50
rect 3434 16 3468 50
rect 3502 16 3536 50
rect 3570 16 3604 50
rect 3638 16 3672 50
rect 3706 16 3740 50
rect 3774 16 3808 50
rect 3842 16 3876 50
rect 3910 16 3944 50
rect 3978 16 4012 50
rect 4046 16 4080 50
rect 4114 16 4148 50
rect 4182 16 4216 50
rect 4250 16 4284 50
rect 4318 16 4352 50
rect 4386 16 4420 50
rect 4454 16 4488 50
rect 4522 16 4556 50
rect 4590 16 4624 50
rect 4658 16 4692 50
rect 4726 16 4760 50
rect 4794 16 4828 50
rect 4862 16 4896 50
rect 4930 16 4964 50
rect 4998 16 5032 50
rect 5066 16 5100 50
rect 5134 16 5168 50
rect 5202 16 5236 50
rect 5270 16 5304 50
rect 5338 16 5372 50
rect 5406 16 5440 50
rect 5474 16 5508 50
rect 5542 16 5576 50
rect 5610 16 5644 50
rect 5678 16 5712 50
rect 5746 16 5780 50
rect 5814 16 5848 50
rect 5882 16 5916 50
rect 5950 16 5984 50
rect 6018 16 6052 50
rect 6086 16 6120 50
rect 6154 16 6188 50
rect 6222 16 6256 50
rect 6290 16 6324 50
rect 6358 16 6392 50
rect 6426 16 6460 50
rect 6494 16 6528 50
rect 6562 16 6596 50
rect 6630 16 6664 50
rect 6698 16 6732 50
rect 6766 16 6800 50
rect 6834 16 6868 50
rect 6902 16 6936 50
rect 6970 16 7004 50
rect 7038 16 7072 50
rect 7106 16 7140 50
rect 7174 16 7208 50
rect 7242 16 7276 50
rect 7310 16 7344 50
rect 7378 16 7412 50
rect 7446 16 7480 50
rect 7514 16 7548 50
rect 7582 16 7616 50
rect 7650 16 7684 50
rect 7718 16 7752 50
rect 7786 16 7820 50
rect 7854 16 7888 50
rect 7922 16 7956 50
rect 7990 16 8024 50
rect 8058 16 8092 50
rect 8126 16 8160 50
rect 8194 16 8228 50
rect 8262 16 8296 50
rect 8330 16 8364 50
rect 8398 16 8432 50
rect 8466 16 8500 50
rect 8534 16 8568 50
rect 8602 16 8636 50
rect 8670 16 8704 50
rect 8738 16 8772 50
rect 8806 16 8840 50
rect 8874 16 8908 50
rect 8942 16 8976 50
rect 9010 16 9044 50
rect 9078 16 9112 50
rect 9146 16 9180 50
rect 9214 16 9248 50
rect 9282 16 9316 50
rect 9350 16 9384 50
rect 9418 16 9452 50
rect 9486 16 9520 50
rect 9554 16 9588 50
rect 9622 16 9656 50
rect 9690 16 9724 50
rect 9758 16 9792 50
rect 9826 16 9860 50
rect 9894 16 9928 50
rect 9962 16 9996 50
rect 10030 16 10064 50
rect 10098 16 10132 50
rect 10166 16 10200 50
rect 10234 16 10268 50
rect 10302 16 10336 50
rect 10370 16 10404 50
rect 10438 16 10472 50
rect 10506 16 10540 50
rect 10574 16 10608 50
rect 10642 16 10676 50
rect 10710 16 10744 50
rect 10778 16 10812 50
rect 10846 16 10880 50
rect 10914 16 10948 50
rect 10982 16 11016 50
rect 11050 16 11084 50
<< locali >>
rect 0 2322 11146 2338
rect 0 2288 34 2322
rect 72 2288 102 2322
rect 144 2288 170 2322
rect 216 2288 238 2322
rect 288 2288 306 2322
rect 360 2288 374 2322
rect 432 2288 442 2322
rect 504 2288 510 2322
rect 576 2288 578 2322
rect 612 2288 614 2322
rect 680 2288 686 2322
rect 748 2288 758 2322
rect 816 2288 830 2322
rect 884 2288 902 2322
rect 952 2288 974 2322
rect 1020 2288 1046 2322
rect 1088 2288 1118 2322
rect 1156 2288 1190 2322
rect 1224 2288 1258 2322
rect 1296 2288 1326 2322
rect 1368 2288 1394 2322
rect 1440 2288 1462 2322
rect 1512 2288 1530 2322
rect 1584 2288 1598 2322
rect 1656 2288 1666 2322
rect 1728 2288 1734 2322
rect 1800 2288 1802 2322
rect 1836 2288 1838 2322
rect 1904 2288 1910 2322
rect 1972 2288 1982 2322
rect 2040 2288 2054 2322
rect 2108 2288 2126 2322
rect 2176 2288 2198 2322
rect 2244 2288 2270 2322
rect 2312 2288 2342 2322
rect 2380 2288 2414 2322
rect 2448 2288 2482 2322
rect 2520 2288 2550 2322
rect 2592 2288 2618 2322
rect 2664 2288 2686 2322
rect 2736 2288 2754 2322
rect 2808 2288 2822 2322
rect 2880 2288 2890 2322
rect 2952 2288 2958 2322
rect 3024 2288 3026 2322
rect 3060 2288 3062 2322
rect 3128 2288 3134 2322
rect 3196 2288 3206 2322
rect 3264 2288 3278 2322
rect 3332 2288 3350 2322
rect 3400 2288 3422 2322
rect 3468 2288 3494 2322
rect 3536 2288 3566 2322
rect 3604 2288 3638 2322
rect 3672 2288 3706 2322
rect 3744 2288 3774 2322
rect 3816 2288 3842 2322
rect 3888 2288 3910 2322
rect 3960 2288 3978 2322
rect 4032 2288 4046 2322
rect 4104 2288 4114 2322
rect 4176 2288 4182 2322
rect 4248 2288 4250 2322
rect 4284 2288 4286 2322
rect 4352 2288 4358 2322
rect 4420 2288 4430 2322
rect 4488 2288 4502 2322
rect 4556 2288 4574 2322
rect 4624 2288 4646 2322
rect 4692 2288 4718 2322
rect 4760 2288 4790 2322
rect 4828 2288 4862 2322
rect 4896 2288 4930 2322
rect 4968 2288 4998 2322
rect 5040 2288 5066 2322
rect 5112 2288 5134 2322
rect 5184 2288 5202 2322
rect 5256 2288 5270 2322
rect 5328 2288 5338 2322
rect 5400 2288 5406 2322
rect 5472 2288 5474 2322
rect 5508 2288 5510 2322
rect 5576 2288 5582 2322
rect 5644 2288 5654 2322
rect 5712 2288 5726 2322
rect 5780 2288 5798 2322
rect 5848 2288 5870 2322
rect 5916 2288 5942 2322
rect 5984 2288 6014 2322
rect 6052 2288 6086 2322
rect 6120 2288 6154 2322
rect 6192 2288 6222 2322
rect 6264 2288 6290 2322
rect 6336 2288 6358 2322
rect 6408 2288 6426 2322
rect 6480 2288 6494 2322
rect 6552 2288 6562 2322
rect 6624 2288 6630 2322
rect 6696 2288 6698 2322
rect 6732 2288 6734 2322
rect 6800 2288 6806 2322
rect 6868 2288 6878 2322
rect 6936 2288 6950 2322
rect 7004 2288 7022 2322
rect 7072 2288 7094 2322
rect 7140 2288 7166 2322
rect 7208 2288 7238 2322
rect 7276 2288 7310 2322
rect 7344 2288 7378 2322
rect 7416 2288 7446 2322
rect 7488 2288 7514 2322
rect 7560 2288 7582 2322
rect 7632 2288 7650 2322
rect 7704 2288 7718 2322
rect 7776 2288 7786 2322
rect 7848 2288 7854 2322
rect 7920 2288 7922 2322
rect 7956 2288 7958 2322
rect 8024 2288 8030 2322
rect 8092 2288 8102 2322
rect 8160 2288 8174 2322
rect 8228 2288 8246 2322
rect 8296 2288 8318 2322
rect 8364 2288 8390 2322
rect 8432 2288 8462 2322
rect 8500 2288 8534 2322
rect 8568 2288 8602 2322
rect 8640 2288 8670 2322
rect 8712 2288 8738 2322
rect 8784 2288 8806 2322
rect 8856 2288 8874 2322
rect 8928 2288 8942 2322
rect 9000 2288 9010 2322
rect 9072 2288 9078 2322
rect 9144 2288 9146 2322
rect 9180 2288 9182 2322
rect 9248 2288 9254 2322
rect 9316 2288 9326 2322
rect 9384 2288 9398 2322
rect 9452 2288 9470 2322
rect 9520 2288 9542 2322
rect 9588 2288 9614 2322
rect 9656 2288 9686 2322
rect 9724 2288 9758 2322
rect 9792 2288 9826 2322
rect 9864 2288 9894 2322
rect 9936 2288 9962 2322
rect 10008 2288 10030 2322
rect 10080 2288 10098 2322
rect 10152 2288 10166 2322
rect 10224 2288 10234 2322
rect 10296 2288 10302 2322
rect 10368 2288 10370 2322
rect 10404 2288 10406 2322
rect 10472 2288 10478 2322
rect 10540 2288 10550 2322
rect 10608 2288 10622 2322
rect 10676 2288 10694 2322
rect 10744 2288 10766 2322
rect 10812 2288 10838 2322
rect 10880 2288 10910 2322
rect 10948 2288 10982 2322
rect 11016 2288 11050 2322
rect 11088 2288 11146 2322
rect 0 2272 11146 2288
rect 0 66 28 2244
rect 56 94 84 2272
rect 112 66 140 2244
rect 168 94 196 2272
rect 224 66 252 2244
rect 280 94 308 2272
rect 336 66 364 2244
rect 392 94 420 2272
rect 448 66 476 2244
rect 504 94 532 2272
rect 560 66 588 2244
rect 616 94 644 2272
rect 672 66 700 2244
rect 728 94 756 2272
rect 784 66 812 2244
rect 840 94 868 2272
rect 896 66 924 2244
rect 952 94 980 2272
rect 1008 66 1036 2244
rect 1064 94 1092 2272
rect 1120 66 1148 2244
rect 1176 94 1204 2272
rect 1232 66 1260 2244
rect 1288 94 1316 2272
rect 1344 66 1372 2244
rect 1400 94 1428 2272
rect 1456 66 1484 2244
rect 1512 94 1540 2272
rect 1568 66 1596 2244
rect 1624 94 1652 2272
rect 1680 66 1708 2244
rect 1736 94 1764 2272
rect 1792 66 1820 2244
rect 1848 94 1876 2272
rect 1904 66 1932 2244
rect 1960 94 1988 2272
rect 2016 66 2044 2244
rect 2072 94 2100 2272
rect 2128 66 2156 2244
rect 2184 94 2212 2272
rect 2240 66 2268 2244
rect 2296 94 2324 2272
rect 2352 66 2380 2244
rect 2408 94 2436 2272
rect 2464 66 2492 2244
rect 2520 94 2548 2272
rect 2576 66 2604 2244
rect 2632 94 2660 2272
rect 2688 66 2716 2244
rect 2744 94 2772 2272
rect 2800 66 2828 2244
rect 2856 94 2884 2272
rect 2912 66 2940 2244
rect 2968 94 2996 2272
rect 3024 66 3052 2244
rect 3080 94 3108 2272
rect 3136 66 3164 2244
rect 3192 94 3220 2272
rect 3248 66 3276 2244
rect 3304 94 3332 2272
rect 3360 66 3388 2244
rect 3416 94 3444 2272
rect 3472 66 3500 2244
rect 3528 94 3556 2272
rect 3584 66 3612 2244
rect 3640 94 3668 2272
rect 3696 66 3724 2244
rect 3752 94 3780 2272
rect 3808 66 3836 2244
rect 3864 94 3892 2272
rect 3920 66 3948 2244
rect 3976 94 4004 2272
rect 4032 66 4060 2244
rect 4088 94 4116 2272
rect 4144 66 4172 2244
rect 4200 94 4228 2272
rect 4256 66 4284 2244
rect 4312 94 4340 2272
rect 4368 66 4396 2244
rect 4424 94 4452 2272
rect 4480 66 4508 2244
rect 4536 94 4564 2272
rect 4592 66 4620 2244
rect 4648 94 4676 2272
rect 4704 66 4732 2244
rect 4760 94 4788 2272
rect 4816 66 4844 2244
rect 4872 94 4900 2272
rect 4928 66 4956 2244
rect 4984 94 5012 2272
rect 5040 66 5068 2244
rect 5096 94 5124 2272
rect 5152 66 5180 2244
rect 5208 94 5236 2272
rect 5264 66 5292 2244
rect 5320 94 5348 2272
rect 5376 66 5404 2244
rect 5432 94 5460 2272
rect 5488 66 5516 2244
rect 5544 94 5572 2272
rect 5600 66 5628 2244
rect 5656 94 5684 2272
rect 5712 66 5740 2244
rect 5768 94 5796 2272
rect 5824 66 5852 2244
rect 5880 94 5908 2272
rect 5936 66 5964 2244
rect 5992 94 6020 2272
rect 6048 66 6076 2244
rect 6104 94 6132 2272
rect 6160 66 6188 2244
rect 6216 94 6244 2272
rect 6272 66 6300 2244
rect 6328 94 6356 2272
rect 6384 66 6412 2244
rect 6440 94 6468 2272
rect 6496 66 6524 2244
rect 6552 94 6580 2272
rect 6608 66 6636 2244
rect 6664 94 6692 2272
rect 6720 66 6748 2244
rect 6776 94 6804 2272
rect 6832 66 6860 2244
rect 6888 94 6916 2272
rect 6944 66 6972 2244
rect 7000 94 7028 2272
rect 7056 66 7084 2244
rect 7112 94 7140 2272
rect 7168 66 7196 2244
rect 7224 94 7252 2272
rect 7280 66 7308 2244
rect 7336 94 7364 2272
rect 7392 66 7420 2244
rect 7448 94 7476 2272
rect 7504 66 7532 2244
rect 7560 94 7588 2272
rect 7616 66 7644 2244
rect 7672 94 7700 2272
rect 7728 66 7756 2244
rect 7784 94 7812 2272
rect 7840 66 7868 2244
rect 7896 94 7924 2272
rect 7952 66 7980 2244
rect 8008 94 8036 2272
rect 8064 66 8092 2244
rect 8120 94 8148 2272
rect 8176 66 8204 2244
rect 8232 94 8260 2272
rect 8288 66 8316 2244
rect 8344 94 8372 2272
rect 8400 66 8428 2244
rect 8456 94 8484 2272
rect 8512 66 8540 2244
rect 8568 94 8596 2272
rect 8624 66 8652 2244
rect 8680 94 8708 2272
rect 8736 66 8764 2244
rect 8792 94 8820 2272
rect 8848 66 8876 2244
rect 8904 94 8932 2272
rect 8960 66 8988 2244
rect 9016 94 9044 2272
rect 9072 66 9100 2244
rect 9128 94 9156 2272
rect 9184 66 9212 2244
rect 9240 94 9268 2272
rect 9296 66 9324 2244
rect 9352 94 9380 2272
rect 9408 66 9436 2244
rect 9464 94 9492 2272
rect 9520 66 9548 2244
rect 9576 94 9604 2272
rect 9632 66 9660 2244
rect 9688 94 9716 2272
rect 9744 66 9772 2244
rect 9800 94 9828 2272
rect 9856 66 9884 2244
rect 9912 94 9940 2272
rect 9968 66 9996 2244
rect 10024 94 10052 2272
rect 10080 66 10108 2244
rect 10136 94 10164 2272
rect 10192 66 10220 2244
rect 10248 94 10276 2272
rect 10304 66 10332 2244
rect 10360 94 10388 2272
rect 10416 66 10444 2244
rect 10472 94 10500 2272
rect 10528 66 10556 2244
rect 10584 94 10612 2272
rect 10640 66 10668 2244
rect 10696 94 10724 2272
rect 10752 66 10780 2244
rect 10808 94 10836 2272
rect 10864 66 10892 2244
rect 10920 94 10948 2272
rect 10976 66 11004 2244
rect 11032 94 11060 2272
rect 11088 66 11146 2244
rect 0 50 11146 66
rect 0 16 34 50
rect 72 16 102 50
rect 144 16 170 50
rect 216 16 238 50
rect 288 16 306 50
rect 360 16 374 50
rect 432 16 442 50
rect 504 16 510 50
rect 576 16 578 50
rect 612 16 614 50
rect 680 16 686 50
rect 748 16 758 50
rect 816 16 830 50
rect 884 16 902 50
rect 952 16 974 50
rect 1020 16 1046 50
rect 1088 16 1118 50
rect 1156 16 1190 50
rect 1224 16 1258 50
rect 1296 16 1326 50
rect 1368 16 1394 50
rect 1440 16 1462 50
rect 1512 16 1530 50
rect 1584 16 1598 50
rect 1656 16 1666 50
rect 1728 16 1734 50
rect 1800 16 1802 50
rect 1836 16 1838 50
rect 1904 16 1910 50
rect 1972 16 1982 50
rect 2040 16 2054 50
rect 2108 16 2126 50
rect 2176 16 2198 50
rect 2244 16 2270 50
rect 2312 16 2342 50
rect 2380 16 2414 50
rect 2448 16 2482 50
rect 2520 16 2550 50
rect 2592 16 2618 50
rect 2664 16 2686 50
rect 2736 16 2754 50
rect 2808 16 2822 50
rect 2880 16 2890 50
rect 2952 16 2958 50
rect 3024 16 3026 50
rect 3060 16 3062 50
rect 3128 16 3134 50
rect 3196 16 3206 50
rect 3264 16 3278 50
rect 3332 16 3350 50
rect 3400 16 3422 50
rect 3468 16 3494 50
rect 3536 16 3566 50
rect 3604 16 3638 50
rect 3672 16 3706 50
rect 3744 16 3774 50
rect 3816 16 3842 50
rect 3888 16 3910 50
rect 3960 16 3978 50
rect 4032 16 4046 50
rect 4104 16 4114 50
rect 4176 16 4182 50
rect 4248 16 4250 50
rect 4284 16 4286 50
rect 4352 16 4358 50
rect 4420 16 4430 50
rect 4488 16 4502 50
rect 4556 16 4574 50
rect 4624 16 4646 50
rect 4692 16 4718 50
rect 4760 16 4790 50
rect 4828 16 4862 50
rect 4896 16 4930 50
rect 4968 16 4998 50
rect 5040 16 5066 50
rect 5112 16 5134 50
rect 5184 16 5202 50
rect 5256 16 5270 50
rect 5328 16 5338 50
rect 5400 16 5406 50
rect 5472 16 5474 50
rect 5508 16 5510 50
rect 5576 16 5582 50
rect 5644 16 5654 50
rect 5712 16 5726 50
rect 5780 16 5798 50
rect 5848 16 5870 50
rect 5916 16 5942 50
rect 5984 16 6014 50
rect 6052 16 6086 50
rect 6120 16 6154 50
rect 6192 16 6222 50
rect 6264 16 6290 50
rect 6336 16 6358 50
rect 6408 16 6426 50
rect 6480 16 6494 50
rect 6552 16 6562 50
rect 6624 16 6630 50
rect 6696 16 6698 50
rect 6732 16 6734 50
rect 6800 16 6806 50
rect 6868 16 6878 50
rect 6936 16 6950 50
rect 7004 16 7022 50
rect 7072 16 7094 50
rect 7140 16 7166 50
rect 7208 16 7238 50
rect 7276 16 7310 50
rect 7344 16 7378 50
rect 7416 16 7446 50
rect 7488 16 7514 50
rect 7560 16 7582 50
rect 7632 16 7650 50
rect 7704 16 7718 50
rect 7776 16 7786 50
rect 7848 16 7854 50
rect 7920 16 7922 50
rect 7956 16 7958 50
rect 8024 16 8030 50
rect 8092 16 8102 50
rect 8160 16 8174 50
rect 8228 16 8246 50
rect 8296 16 8318 50
rect 8364 16 8390 50
rect 8432 16 8462 50
rect 8500 16 8534 50
rect 8568 16 8602 50
rect 8640 16 8670 50
rect 8712 16 8738 50
rect 8784 16 8806 50
rect 8856 16 8874 50
rect 8928 16 8942 50
rect 9000 16 9010 50
rect 9072 16 9078 50
rect 9144 16 9146 50
rect 9180 16 9182 50
rect 9248 16 9254 50
rect 9316 16 9326 50
rect 9384 16 9398 50
rect 9452 16 9470 50
rect 9520 16 9542 50
rect 9588 16 9614 50
rect 9656 16 9686 50
rect 9724 16 9758 50
rect 9792 16 9826 50
rect 9864 16 9894 50
rect 9936 16 9962 50
rect 10008 16 10030 50
rect 10080 16 10098 50
rect 10152 16 10166 50
rect 10224 16 10234 50
rect 10296 16 10302 50
rect 10368 16 10370 50
rect 10404 16 10406 50
rect 10472 16 10478 50
rect 10540 16 10550 50
rect 10608 16 10622 50
rect 10676 16 10694 50
rect 10744 16 10766 50
rect 10812 16 10838 50
rect 10880 16 10910 50
rect 10948 16 10982 50
rect 11016 16 11050 50
rect 11088 16 11146 50
rect 0 0 11146 16
<< viali >>
rect 38 2288 68 2322
rect 68 2288 72 2322
rect 110 2288 136 2322
rect 136 2288 144 2322
rect 182 2288 204 2322
rect 204 2288 216 2322
rect 254 2288 272 2322
rect 272 2288 288 2322
rect 326 2288 340 2322
rect 340 2288 360 2322
rect 398 2288 408 2322
rect 408 2288 432 2322
rect 470 2288 476 2322
rect 476 2288 504 2322
rect 542 2288 544 2322
rect 544 2288 576 2322
rect 614 2288 646 2322
rect 646 2288 648 2322
rect 686 2288 714 2322
rect 714 2288 720 2322
rect 758 2288 782 2322
rect 782 2288 792 2322
rect 830 2288 850 2322
rect 850 2288 864 2322
rect 902 2288 918 2322
rect 918 2288 936 2322
rect 974 2288 986 2322
rect 986 2288 1008 2322
rect 1046 2288 1054 2322
rect 1054 2288 1080 2322
rect 1118 2288 1122 2322
rect 1122 2288 1152 2322
rect 1190 2288 1224 2322
rect 1262 2288 1292 2322
rect 1292 2288 1296 2322
rect 1334 2288 1360 2322
rect 1360 2288 1368 2322
rect 1406 2288 1428 2322
rect 1428 2288 1440 2322
rect 1478 2288 1496 2322
rect 1496 2288 1512 2322
rect 1550 2288 1564 2322
rect 1564 2288 1584 2322
rect 1622 2288 1632 2322
rect 1632 2288 1656 2322
rect 1694 2288 1700 2322
rect 1700 2288 1728 2322
rect 1766 2288 1768 2322
rect 1768 2288 1800 2322
rect 1838 2288 1870 2322
rect 1870 2288 1872 2322
rect 1910 2288 1938 2322
rect 1938 2288 1944 2322
rect 1982 2288 2006 2322
rect 2006 2288 2016 2322
rect 2054 2288 2074 2322
rect 2074 2288 2088 2322
rect 2126 2288 2142 2322
rect 2142 2288 2160 2322
rect 2198 2288 2210 2322
rect 2210 2288 2232 2322
rect 2270 2288 2278 2322
rect 2278 2288 2304 2322
rect 2342 2288 2346 2322
rect 2346 2288 2376 2322
rect 2414 2288 2448 2322
rect 2486 2288 2516 2322
rect 2516 2288 2520 2322
rect 2558 2288 2584 2322
rect 2584 2288 2592 2322
rect 2630 2288 2652 2322
rect 2652 2288 2664 2322
rect 2702 2288 2720 2322
rect 2720 2288 2736 2322
rect 2774 2288 2788 2322
rect 2788 2288 2808 2322
rect 2846 2288 2856 2322
rect 2856 2288 2880 2322
rect 2918 2288 2924 2322
rect 2924 2288 2952 2322
rect 2990 2288 2992 2322
rect 2992 2288 3024 2322
rect 3062 2288 3094 2322
rect 3094 2288 3096 2322
rect 3134 2288 3162 2322
rect 3162 2288 3168 2322
rect 3206 2288 3230 2322
rect 3230 2288 3240 2322
rect 3278 2288 3298 2322
rect 3298 2288 3312 2322
rect 3350 2288 3366 2322
rect 3366 2288 3384 2322
rect 3422 2288 3434 2322
rect 3434 2288 3456 2322
rect 3494 2288 3502 2322
rect 3502 2288 3528 2322
rect 3566 2288 3570 2322
rect 3570 2288 3600 2322
rect 3638 2288 3672 2322
rect 3710 2288 3740 2322
rect 3740 2288 3744 2322
rect 3782 2288 3808 2322
rect 3808 2288 3816 2322
rect 3854 2288 3876 2322
rect 3876 2288 3888 2322
rect 3926 2288 3944 2322
rect 3944 2288 3960 2322
rect 3998 2288 4012 2322
rect 4012 2288 4032 2322
rect 4070 2288 4080 2322
rect 4080 2288 4104 2322
rect 4142 2288 4148 2322
rect 4148 2288 4176 2322
rect 4214 2288 4216 2322
rect 4216 2288 4248 2322
rect 4286 2288 4318 2322
rect 4318 2288 4320 2322
rect 4358 2288 4386 2322
rect 4386 2288 4392 2322
rect 4430 2288 4454 2322
rect 4454 2288 4464 2322
rect 4502 2288 4522 2322
rect 4522 2288 4536 2322
rect 4574 2288 4590 2322
rect 4590 2288 4608 2322
rect 4646 2288 4658 2322
rect 4658 2288 4680 2322
rect 4718 2288 4726 2322
rect 4726 2288 4752 2322
rect 4790 2288 4794 2322
rect 4794 2288 4824 2322
rect 4862 2288 4896 2322
rect 4934 2288 4964 2322
rect 4964 2288 4968 2322
rect 5006 2288 5032 2322
rect 5032 2288 5040 2322
rect 5078 2288 5100 2322
rect 5100 2288 5112 2322
rect 5150 2288 5168 2322
rect 5168 2288 5184 2322
rect 5222 2288 5236 2322
rect 5236 2288 5256 2322
rect 5294 2288 5304 2322
rect 5304 2288 5328 2322
rect 5366 2288 5372 2322
rect 5372 2288 5400 2322
rect 5438 2288 5440 2322
rect 5440 2288 5472 2322
rect 5510 2288 5542 2322
rect 5542 2288 5544 2322
rect 5582 2288 5610 2322
rect 5610 2288 5616 2322
rect 5654 2288 5678 2322
rect 5678 2288 5688 2322
rect 5726 2288 5746 2322
rect 5746 2288 5760 2322
rect 5798 2288 5814 2322
rect 5814 2288 5832 2322
rect 5870 2288 5882 2322
rect 5882 2288 5904 2322
rect 5942 2288 5950 2322
rect 5950 2288 5976 2322
rect 6014 2288 6018 2322
rect 6018 2288 6048 2322
rect 6086 2288 6120 2322
rect 6158 2288 6188 2322
rect 6188 2288 6192 2322
rect 6230 2288 6256 2322
rect 6256 2288 6264 2322
rect 6302 2288 6324 2322
rect 6324 2288 6336 2322
rect 6374 2288 6392 2322
rect 6392 2288 6408 2322
rect 6446 2288 6460 2322
rect 6460 2288 6480 2322
rect 6518 2288 6528 2322
rect 6528 2288 6552 2322
rect 6590 2288 6596 2322
rect 6596 2288 6624 2322
rect 6662 2288 6664 2322
rect 6664 2288 6696 2322
rect 6734 2288 6766 2322
rect 6766 2288 6768 2322
rect 6806 2288 6834 2322
rect 6834 2288 6840 2322
rect 6878 2288 6902 2322
rect 6902 2288 6912 2322
rect 6950 2288 6970 2322
rect 6970 2288 6984 2322
rect 7022 2288 7038 2322
rect 7038 2288 7056 2322
rect 7094 2288 7106 2322
rect 7106 2288 7128 2322
rect 7166 2288 7174 2322
rect 7174 2288 7200 2322
rect 7238 2288 7242 2322
rect 7242 2288 7272 2322
rect 7310 2288 7344 2322
rect 7382 2288 7412 2322
rect 7412 2288 7416 2322
rect 7454 2288 7480 2322
rect 7480 2288 7488 2322
rect 7526 2288 7548 2322
rect 7548 2288 7560 2322
rect 7598 2288 7616 2322
rect 7616 2288 7632 2322
rect 7670 2288 7684 2322
rect 7684 2288 7704 2322
rect 7742 2288 7752 2322
rect 7752 2288 7776 2322
rect 7814 2288 7820 2322
rect 7820 2288 7848 2322
rect 7886 2288 7888 2322
rect 7888 2288 7920 2322
rect 7958 2288 7990 2322
rect 7990 2288 7992 2322
rect 8030 2288 8058 2322
rect 8058 2288 8064 2322
rect 8102 2288 8126 2322
rect 8126 2288 8136 2322
rect 8174 2288 8194 2322
rect 8194 2288 8208 2322
rect 8246 2288 8262 2322
rect 8262 2288 8280 2322
rect 8318 2288 8330 2322
rect 8330 2288 8352 2322
rect 8390 2288 8398 2322
rect 8398 2288 8424 2322
rect 8462 2288 8466 2322
rect 8466 2288 8496 2322
rect 8534 2288 8568 2322
rect 8606 2288 8636 2322
rect 8636 2288 8640 2322
rect 8678 2288 8704 2322
rect 8704 2288 8712 2322
rect 8750 2288 8772 2322
rect 8772 2288 8784 2322
rect 8822 2288 8840 2322
rect 8840 2288 8856 2322
rect 8894 2288 8908 2322
rect 8908 2288 8928 2322
rect 8966 2288 8976 2322
rect 8976 2288 9000 2322
rect 9038 2288 9044 2322
rect 9044 2288 9072 2322
rect 9110 2288 9112 2322
rect 9112 2288 9144 2322
rect 9182 2288 9214 2322
rect 9214 2288 9216 2322
rect 9254 2288 9282 2322
rect 9282 2288 9288 2322
rect 9326 2288 9350 2322
rect 9350 2288 9360 2322
rect 9398 2288 9418 2322
rect 9418 2288 9432 2322
rect 9470 2288 9486 2322
rect 9486 2288 9504 2322
rect 9542 2288 9554 2322
rect 9554 2288 9576 2322
rect 9614 2288 9622 2322
rect 9622 2288 9648 2322
rect 9686 2288 9690 2322
rect 9690 2288 9720 2322
rect 9758 2288 9792 2322
rect 9830 2288 9860 2322
rect 9860 2288 9864 2322
rect 9902 2288 9928 2322
rect 9928 2288 9936 2322
rect 9974 2288 9996 2322
rect 9996 2288 10008 2322
rect 10046 2288 10064 2322
rect 10064 2288 10080 2322
rect 10118 2288 10132 2322
rect 10132 2288 10152 2322
rect 10190 2288 10200 2322
rect 10200 2288 10224 2322
rect 10262 2288 10268 2322
rect 10268 2288 10296 2322
rect 10334 2288 10336 2322
rect 10336 2288 10368 2322
rect 10406 2288 10438 2322
rect 10438 2288 10440 2322
rect 10478 2288 10506 2322
rect 10506 2288 10512 2322
rect 10550 2288 10574 2322
rect 10574 2288 10584 2322
rect 10622 2288 10642 2322
rect 10642 2288 10656 2322
rect 10694 2288 10710 2322
rect 10710 2288 10728 2322
rect 10766 2288 10778 2322
rect 10778 2288 10800 2322
rect 10838 2288 10846 2322
rect 10846 2288 10872 2322
rect 10910 2288 10914 2322
rect 10914 2288 10944 2322
rect 10982 2288 11016 2322
rect 11054 2288 11084 2322
rect 11084 2288 11088 2322
rect 38 16 68 50
rect 68 16 72 50
rect 110 16 136 50
rect 136 16 144 50
rect 182 16 204 50
rect 204 16 216 50
rect 254 16 272 50
rect 272 16 288 50
rect 326 16 340 50
rect 340 16 360 50
rect 398 16 408 50
rect 408 16 432 50
rect 470 16 476 50
rect 476 16 504 50
rect 542 16 544 50
rect 544 16 576 50
rect 614 16 646 50
rect 646 16 648 50
rect 686 16 714 50
rect 714 16 720 50
rect 758 16 782 50
rect 782 16 792 50
rect 830 16 850 50
rect 850 16 864 50
rect 902 16 918 50
rect 918 16 936 50
rect 974 16 986 50
rect 986 16 1008 50
rect 1046 16 1054 50
rect 1054 16 1080 50
rect 1118 16 1122 50
rect 1122 16 1152 50
rect 1190 16 1224 50
rect 1262 16 1292 50
rect 1292 16 1296 50
rect 1334 16 1360 50
rect 1360 16 1368 50
rect 1406 16 1428 50
rect 1428 16 1440 50
rect 1478 16 1496 50
rect 1496 16 1512 50
rect 1550 16 1564 50
rect 1564 16 1584 50
rect 1622 16 1632 50
rect 1632 16 1656 50
rect 1694 16 1700 50
rect 1700 16 1728 50
rect 1766 16 1768 50
rect 1768 16 1800 50
rect 1838 16 1870 50
rect 1870 16 1872 50
rect 1910 16 1938 50
rect 1938 16 1944 50
rect 1982 16 2006 50
rect 2006 16 2016 50
rect 2054 16 2074 50
rect 2074 16 2088 50
rect 2126 16 2142 50
rect 2142 16 2160 50
rect 2198 16 2210 50
rect 2210 16 2232 50
rect 2270 16 2278 50
rect 2278 16 2304 50
rect 2342 16 2346 50
rect 2346 16 2376 50
rect 2414 16 2448 50
rect 2486 16 2516 50
rect 2516 16 2520 50
rect 2558 16 2584 50
rect 2584 16 2592 50
rect 2630 16 2652 50
rect 2652 16 2664 50
rect 2702 16 2720 50
rect 2720 16 2736 50
rect 2774 16 2788 50
rect 2788 16 2808 50
rect 2846 16 2856 50
rect 2856 16 2880 50
rect 2918 16 2924 50
rect 2924 16 2952 50
rect 2990 16 2992 50
rect 2992 16 3024 50
rect 3062 16 3094 50
rect 3094 16 3096 50
rect 3134 16 3162 50
rect 3162 16 3168 50
rect 3206 16 3230 50
rect 3230 16 3240 50
rect 3278 16 3298 50
rect 3298 16 3312 50
rect 3350 16 3366 50
rect 3366 16 3384 50
rect 3422 16 3434 50
rect 3434 16 3456 50
rect 3494 16 3502 50
rect 3502 16 3528 50
rect 3566 16 3570 50
rect 3570 16 3600 50
rect 3638 16 3672 50
rect 3710 16 3740 50
rect 3740 16 3744 50
rect 3782 16 3808 50
rect 3808 16 3816 50
rect 3854 16 3876 50
rect 3876 16 3888 50
rect 3926 16 3944 50
rect 3944 16 3960 50
rect 3998 16 4012 50
rect 4012 16 4032 50
rect 4070 16 4080 50
rect 4080 16 4104 50
rect 4142 16 4148 50
rect 4148 16 4176 50
rect 4214 16 4216 50
rect 4216 16 4248 50
rect 4286 16 4318 50
rect 4318 16 4320 50
rect 4358 16 4386 50
rect 4386 16 4392 50
rect 4430 16 4454 50
rect 4454 16 4464 50
rect 4502 16 4522 50
rect 4522 16 4536 50
rect 4574 16 4590 50
rect 4590 16 4608 50
rect 4646 16 4658 50
rect 4658 16 4680 50
rect 4718 16 4726 50
rect 4726 16 4752 50
rect 4790 16 4794 50
rect 4794 16 4824 50
rect 4862 16 4896 50
rect 4934 16 4964 50
rect 4964 16 4968 50
rect 5006 16 5032 50
rect 5032 16 5040 50
rect 5078 16 5100 50
rect 5100 16 5112 50
rect 5150 16 5168 50
rect 5168 16 5184 50
rect 5222 16 5236 50
rect 5236 16 5256 50
rect 5294 16 5304 50
rect 5304 16 5328 50
rect 5366 16 5372 50
rect 5372 16 5400 50
rect 5438 16 5440 50
rect 5440 16 5472 50
rect 5510 16 5542 50
rect 5542 16 5544 50
rect 5582 16 5610 50
rect 5610 16 5616 50
rect 5654 16 5678 50
rect 5678 16 5688 50
rect 5726 16 5746 50
rect 5746 16 5760 50
rect 5798 16 5814 50
rect 5814 16 5832 50
rect 5870 16 5882 50
rect 5882 16 5904 50
rect 5942 16 5950 50
rect 5950 16 5976 50
rect 6014 16 6018 50
rect 6018 16 6048 50
rect 6086 16 6120 50
rect 6158 16 6188 50
rect 6188 16 6192 50
rect 6230 16 6256 50
rect 6256 16 6264 50
rect 6302 16 6324 50
rect 6324 16 6336 50
rect 6374 16 6392 50
rect 6392 16 6408 50
rect 6446 16 6460 50
rect 6460 16 6480 50
rect 6518 16 6528 50
rect 6528 16 6552 50
rect 6590 16 6596 50
rect 6596 16 6624 50
rect 6662 16 6664 50
rect 6664 16 6696 50
rect 6734 16 6766 50
rect 6766 16 6768 50
rect 6806 16 6834 50
rect 6834 16 6840 50
rect 6878 16 6902 50
rect 6902 16 6912 50
rect 6950 16 6970 50
rect 6970 16 6984 50
rect 7022 16 7038 50
rect 7038 16 7056 50
rect 7094 16 7106 50
rect 7106 16 7128 50
rect 7166 16 7174 50
rect 7174 16 7200 50
rect 7238 16 7242 50
rect 7242 16 7272 50
rect 7310 16 7344 50
rect 7382 16 7412 50
rect 7412 16 7416 50
rect 7454 16 7480 50
rect 7480 16 7488 50
rect 7526 16 7548 50
rect 7548 16 7560 50
rect 7598 16 7616 50
rect 7616 16 7632 50
rect 7670 16 7684 50
rect 7684 16 7704 50
rect 7742 16 7752 50
rect 7752 16 7776 50
rect 7814 16 7820 50
rect 7820 16 7848 50
rect 7886 16 7888 50
rect 7888 16 7920 50
rect 7958 16 7990 50
rect 7990 16 7992 50
rect 8030 16 8058 50
rect 8058 16 8064 50
rect 8102 16 8126 50
rect 8126 16 8136 50
rect 8174 16 8194 50
rect 8194 16 8208 50
rect 8246 16 8262 50
rect 8262 16 8280 50
rect 8318 16 8330 50
rect 8330 16 8352 50
rect 8390 16 8398 50
rect 8398 16 8424 50
rect 8462 16 8466 50
rect 8466 16 8496 50
rect 8534 16 8568 50
rect 8606 16 8636 50
rect 8636 16 8640 50
rect 8678 16 8704 50
rect 8704 16 8712 50
rect 8750 16 8772 50
rect 8772 16 8784 50
rect 8822 16 8840 50
rect 8840 16 8856 50
rect 8894 16 8908 50
rect 8908 16 8928 50
rect 8966 16 8976 50
rect 8976 16 9000 50
rect 9038 16 9044 50
rect 9044 16 9072 50
rect 9110 16 9112 50
rect 9112 16 9144 50
rect 9182 16 9214 50
rect 9214 16 9216 50
rect 9254 16 9282 50
rect 9282 16 9288 50
rect 9326 16 9350 50
rect 9350 16 9360 50
rect 9398 16 9418 50
rect 9418 16 9432 50
rect 9470 16 9486 50
rect 9486 16 9504 50
rect 9542 16 9554 50
rect 9554 16 9576 50
rect 9614 16 9622 50
rect 9622 16 9648 50
rect 9686 16 9690 50
rect 9690 16 9720 50
rect 9758 16 9792 50
rect 9830 16 9860 50
rect 9860 16 9864 50
rect 9902 16 9928 50
rect 9928 16 9936 50
rect 9974 16 9996 50
rect 9996 16 10008 50
rect 10046 16 10064 50
rect 10064 16 10080 50
rect 10118 16 10132 50
rect 10132 16 10152 50
rect 10190 16 10200 50
rect 10200 16 10224 50
rect 10262 16 10268 50
rect 10268 16 10296 50
rect 10334 16 10336 50
rect 10336 16 10368 50
rect 10406 16 10438 50
rect 10438 16 10440 50
rect 10478 16 10506 50
rect 10506 16 10512 50
rect 10550 16 10574 50
rect 10574 16 10584 50
rect 10622 16 10642 50
rect 10642 16 10656 50
rect 10694 16 10710 50
rect 10710 16 10728 50
rect 10766 16 10778 50
rect 10778 16 10800 50
rect 10838 16 10846 50
rect 10846 16 10872 50
rect 10910 16 10914 50
rect 10914 16 10944 50
rect 10982 16 11016 50
rect 11054 16 11084 50
rect 11084 16 11088 50
<< metal1 >>
rect 0 2331 11146 2338
rect 0 2322 68 2331
rect 120 2322 132 2331
rect 184 2322 292 2331
rect 344 2322 356 2331
rect 408 2322 516 2331
rect 568 2322 580 2331
rect 632 2322 740 2331
rect 0 2288 38 2322
rect 216 2288 254 2322
rect 288 2288 292 2322
rect 432 2288 470 2322
rect 504 2288 516 2322
rect 576 2288 580 2322
rect 648 2288 686 2322
rect 720 2288 740 2322
rect 0 2279 68 2288
rect 120 2279 132 2288
rect 184 2279 292 2288
rect 344 2279 356 2288
rect 408 2279 516 2288
rect 568 2279 580 2288
rect 632 2279 740 2288
rect 792 2279 804 2331
rect 856 2322 964 2331
rect 864 2288 902 2322
rect 936 2288 964 2322
rect 856 2279 964 2288
rect 1016 2279 1028 2331
rect 1080 2322 1188 2331
rect 1080 2288 1118 2322
rect 1152 2288 1188 2322
rect 1080 2279 1188 2288
rect 1240 2279 1252 2331
rect 1304 2322 1412 2331
rect 1304 2288 1334 2322
rect 1368 2288 1406 2322
rect 1304 2279 1412 2288
rect 1464 2279 1476 2331
rect 1528 2322 1636 2331
rect 1688 2322 1700 2331
rect 1752 2322 1860 2331
rect 1912 2322 1924 2331
rect 1976 2322 2084 2331
rect 2136 2322 2148 2331
rect 2200 2322 2308 2331
rect 2360 2322 2372 2331
rect 2424 2322 2532 2331
rect 2584 2322 2596 2331
rect 2648 2322 2756 2331
rect 1528 2288 1550 2322
rect 1584 2288 1622 2322
rect 1688 2288 1694 2322
rect 1752 2288 1766 2322
rect 1800 2288 1838 2322
rect 1976 2288 1982 2322
rect 2016 2288 2054 2322
rect 2232 2288 2270 2322
rect 2304 2288 2308 2322
rect 2448 2288 2486 2322
rect 2520 2288 2532 2322
rect 2592 2288 2596 2322
rect 2664 2288 2702 2322
rect 2736 2288 2756 2322
rect 1528 2279 1636 2288
rect 1688 2279 1700 2288
rect 1752 2279 1860 2288
rect 1912 2279 1924 2288
rect 1976 2279 2084 2288
rect 2136 2279 2148 2288
rect 2200 2279 2308 2288
rect 2360 2279 2372 2288
rect 2424 2279 2532 2288
rect 2584 2279 2596 2288
rect 2648 2279 2756 2288
rect 2808 2279 2820 2331
rect 2872 2322 2980 2331
rect 2880 2288 2918 2322
rect 2952 2288 2980 2322
rect 2872 2279 2980 2288
rect 3032 2279 3044 2331
rect 3096 2322 3204 2331
rect 3096 2288 3134 2322
rect 3168 2288 3204 2322
rect 3096 2279 3204 2288
rect 3256 2279 3268 2331
rect 3320 2322 3428 2331
rect 3320 2288 3350 2322
rect 3384 2288 3422 2322
rect 3320 2279 3428 2288
rect 3480 2279 3492 2331
rect 3544 2322 3652 2331
rect 3704 2322 3716 2331
rect 3768 2322 3876 2331
rect 3928 2322 3940 2331
rect 3992 2322 4100 2331
rect 4152 2322 4164 2331
rect 4216 2322 4324 2331
rect 4376 2322 4388 2331
rect 4440 2322 4548 2331
rect 4600 2322 4612 2331
rect 4664 2322 4772 2331
rect 3544 2288 3566 2322
rect 3600 2288 3638 2322
rect 3704 2288 3710 2322
rect 3768 2288 3782 2322
rect 3816 2288 3854 2322
rect 3992 2288 3998 2322
rect 4032 2288 4070 2322
rect 4248 2288 4286 2322
rect 4320 2288 4324 2322
rect 4464 2288 4502 2322
rect 4536 2288 4548 2322
rect 4608 2288 4612 2322
rect 4680 2288 4718 2322
rect 4752 2288 4772 2322
rect 3544 2279 3652 2288
rect 3704 2279 3716 2288
rect 3768 2279 3876 2288
rect 3928 2279 3940 2288
rect 3992 2279 4100 2288
rect 4152 2279 4164 2288
rect 4216 2279 4324 2288
rect 4376 2279 4388 2288
rect 4440 2279 4548 2288
rect 4600 2279 4612 2288
rect 4664 2279 4772 2288
rect 4824 2279 4836 2331
rect 4888 2322 4996 2331
rect 4896 2288 4934 2322
rect 4968 2288 4996 2322
rect 4888 2279 4996 2288
rect 5048 2279 5060 2331
rect 5112 2322 5220 2331
rect 5112 2288 5150 2322
rect 5184 2288 5220 2322
rect 5112 2279 5220 2288
rect 5272 2279 5284 2331
rect 5336 2322 5444 2331
rect 5336 2288 5366 2322
rect 5400 2288 5438 2322
rect 5336 2279 5444 2288
rect 5496 2279 5508 2331
rect 5560 2322 5668 2331
rect 5720 2322 5732 2331
rect 5784 2322 5892 2331
rect 5944 2322 5956 2331
rect 6008 2322 6116 2331
rect 6168 2322 6180 2331
rect 6232 2322 6340 2331
rect 6392 2322 6404 2331
rect 6456 2322 6564 2331
rect 6616 2322 6628 2331
rect 6680 2322 6788 2331
rect 5560 2288 5582 2322
rect 5616 2288 5654 2322
rect 5720 2288 5726 2322
rect 5784 2288 5798 2322
rect 5832 2288 5870 2322
rect 6008 2288 6014 2322
rect 6048 2288 6086 2322
rect 6264 2288 6302 2322
rect 6336 2288 6340 2322
rect 6480 2288 6518 2322
rect 6552 2288 6564 2322
rect 6624 2288 6628 2322
rect 6696 2288 6734 2322
rect 6768 2288 6788 2322
rect 5560 2279 5668 2288
rect 5720 2279 5732 2288
rect 5784 2279 5892 2288
rect 5944 2279 5956 2288
rect 6008 2279 6116 2288
rect 6168 2279 6180 2288
rect 6232 2279 6340 2288
rect 6392 2279 6404 2288
rect 6456 2279 6564 2288
rect 6616 2279 6628 2288
rect 6680 2279 6788 2288
rect 6840 2279 6852 2331
rect 6904 2322 7012 2331
rect 6912 2288 6950 2322
rect 6984 2288 7012 2322
rect 6904 2279 7012 2288
rect 7064 2279 7076 2331
rect 7128 2322 7236 2331
rect 7128 2288 7166 2322
rect 7200 2288 7236 2322
rect 7128 2279 7236 2288
rect 7288 2279 7300 2331
rect 7352 2322 7460 2331
rect 7352 2288 7382 2322
rect 7416 2288 7454 2322
rect 7352 2279 7460 2288
rect 7512 2279 7524 2331
rect 7576 2322 7684 2331
rect 7736 2322 7748 2331
rect 7800 2322 7908 2331
rect 7960 2322 7972 2331
rect 8024 2322 8132 2331
rect 8184 2322 8196 2331
rect 8248 2322 8356 2331
rect 8408 2322 8420 2331
rect 8472 2322 8580 2331
rect 8632 2322 8644 2331
rect 8696 2322 8804 2331
rect 7576 2288 7598 2322
rect 7632 2288 7670 2322
rect 7736 2288 7742 2322
rect 7800 2288 7814 2322
rect 7848 2288 7886 2322
rect 8024 2288 8030 2322
rect 8064 2288 8102 2322
rect 8280 2288 8318 2322
rect 8352 2288 8356 2322
rect 8496 2288 8534 2322
rect 8568 2288 8580 2322
rect 8640 2288 8644 2322
rect 8712 2288 8750 2322
rect 8784 2288 8804 2322
rect 7576 2279 7684 2288
rect 7736 2279 7748 2288
rect 7800 2279 7908 2288
rect 7960 2279 7972 2288
rect 8024 2279 8132 2288
rect 8184 2279 8196 2288
rect 8248 2279 8356 2288
rect 8408 2279 8420 2288
rect 8472 2279 8580 2288
rect 8632 2279 8644 2288
rect 8696 2279 8804 2288
rect 8856 2279 8868 2331
rect 8920 2322 9028 2331
rect 8928 2288 8966 2322
rect 9000 2288 9028 2322
rect 8920 2279 9028 2288
rect 9080 2279 9092 2331
rect 9144 2322 9252 2331
rect 9144 2288 9182 2322
rect 9216 2288 9252 2322
rect 9144 2279 9252 2288
rect 9304 2279 9316 2331
rect 9368 2322 9476 2331
rect 9368 2288 9398 2322
rect 9432 2288 9470 2322
rect 9368 2279 9476 2288
rect 9528 2279 9540 2331
rect 9592 2322 9700 2331
rect 9752 2322 9764 2331
rect 9816 2322 9924 2331
rect 9976 2322 9988 2331
rect 10040 2322 10148 2331
rect 10200 2322 10212 2331
rect 10264 2322 10372 2331
rect 10424 2322 10436 2331
rect 10488 2322 10596 2331
rect 10648 2322 10660 2331
rect 10712 2322 10820 2331
rect 9592 2288 9614 2322
rect 9648 2288 9686 2322
rect 9752 2288 9758 2322
rect 9816 2288 9830 2322
rect 9864 2288 9902 2322
rect 10040 2288 10046 2322
rect 10080 2288 10118 2322
rect 10296 2288 10334 2322
rect 10368 2288 10372 2322
rect 10512 2288 10550 2322
rect 10584 2288 10596 2322
rect 10656 2288 10660 2322
rect 10728 2288 10766 2322
rect 10800 2288 10820 2322
rect 9592 2279 9700 2288
rect 9752 2279 9764 2288
rect 9816 2279 9924 2288
rect 9976 2279 9988 2288
rect 10040 2279 10148 2288
rect 10200 2279 10212 2288
rect 10264 2279 10372 2288
rect 10424 2279 10436 2288
rect 10488 2279 10596 2288
rect 10648 2279 10660 2288
rect 10712 2279 10820 2288
rect 10872 2279 10884 2331
rect 10936 2322 11146 2331
rect 10944 2288 10982 2322
rect 11016 2288 11054 2322
rect 11088 2288 11146 2322
rect 10936 2279 11146 2288
rect 0 2272 11146 2279
rect 0 94 28 2272
rect 56 66 84 2244
rect 112 94 140 2272
rect 168 66 196 2244
rect 224 94 252 2272
rect 280 66 308 2244
rect 336 94 364 2272
rect 392 66 420 2244
rect 448 94 476 2272
rect 504 66 532 2244
rect 560 94 588 2272
rect 616 66 644 2244
rect 672 94 700 2272
rect 728 66 756 2244
rect 784 94 812 2272
rect 840 66 868 2244
rect 896 94 924 2272
rect 952 66 980 2244
rect 1008 94 1036 2272
rect 1064 66 1092 2244
rect 1120 94 1148 2272
rect 1176 66 1204 2244
rect 1232 94 1260 2272
rect 1288 66 1316 2244
rect 1344 94 1372 2272
rect 1400 66 1428 2244
rect 1456 94 1484 2272
rect 1512 66 1540 2244
rect 1568 94 1596 2272
rect 1624 66 1652 2244
rect 1680 94 1708 2272
rect 1736 66 1764 2244
rect 1792 94 1820 2272
rect 1848 66 1876 2244
rect 1904 94 1932 2272
rect 1960 66 1988 2244
rect 2016 94 2044 2272
rect 2072 66 2100 2244
rect 2128 94 2156 2272
rect 2184 66 2212 2244
rect 2240 94 2268 2272
rect 2296 66 2324 2244
rect 2352 94 2380 2272
rect 2408 66 2436 2244
rect 2464 94 2492 2272
rect 2520 66 2548 2244
rect 2576 94 2604 2272
rect 2632 66 2660 2244
rect 2688 94 2716 2272
rect 2744 66 2772 2244
rect 2800 94 2828 2272
rect 2856 66 2884 2244
rect 2912 94 2940 2272
rect 2968 66 2996 2244
rect 3024 94 3052 2272
rect 3080 66 3108 2244
rect 3136 94 3164 2272
rect 3192 66 3220 2244
rect 3248 94 3276 2272
rect 3304 66 3332 2244
rect 3360 94 3388 2272
rect 3416 66 3444 2244
rect 3472 94 3500 2272
rect 3528 66 3556 2244
rect 3584 94 3612 2272
rect 3640 66 3668 2244
rect 3696 94 3724 2272
rect 3752 66 3780 2244
rect 3808 94 3836 2272
rect 3864 66 3892 2244
rect 3920 94 3948 2272
rect 3976 66 4004 2244
rect 4032 94 4060 2272
rect 4088 66 4116 2244
rect 4144 94 4172 2272
rect 4200 66 4228 2244
rect 4256 94 4284 2272
rect 4312 66 4340 2244
rect 4368 94 4396 2272
rect 4424 66 4452 2244
rect 4480 94 4508 2272
rect 4536 66 4564 2244
rect 4592 94 4620 2272
rect 4648 66 4676 2244
rect 4704 94 4732 2272
rect 4760 66 4788 2244
rect 4816 94 4844 2272
rect 4872 66 4900 2244
rect 4928 94 4956 2272
rect 4984 66 5012 2244
rect 5040 94 5068 2272
rect 5096 66 5124 2244
rect 5152 94 5180 2272
rect 5208 66 5236 2244
rect 5264 94 5292 2272
rect 5320 66 5348 2244
rect 5376 94 5404 2272
rect 5432 66 5460 2244
rect 5488 94 5516 2272
rect 5544 66 5572 2244
rect 5600 94 5628 2272
rect 5656 66 5684 2244
rect 5712 94 5740 2272
rect 5768 66 5796 2244
rect 5824 94 5852 2272
rect 5880 66 5908 2244
rect 5936 94 5964 2272
rect 5992 66 6020 2244
rect 6048 94 6076 2272
rect 6104 66 6132 2244
rect 6160 94 6188 2272
rect 6216 66 6244 2244
rect 6272 94 6300 2272
rect 6328 66 6356 2244
rect 6384 94 6412 2272
rect 6440 66 6468 2244
rect 6496 94 6524 2272
rect 6552 66 6580 2244
rect 6608 94 6636 2272
rect 6664 66 6692 2244
rect 6720 94 6748 2272
rect 6776 66 6804 2244
rect 6832 94 6860 2272
rect 6888 66 6916 2244
rect 6944 94 6972 2272
rect 7000 66 7028 2244
rect 7056 94 7084 2272
rect 7112 66 7140 2244
rect 7168 94 7196 2272
rect 7224 66 7252 2244
rect 7280 94 7308 2272
rect 7336 66 7364 2244
rect 7392 94 7420 2272
rect 7448 66 7476 2244
rect 7504 94 7532 2272
rect 7560 66 7588 2244
rect 7616 94 7644 2272
rect 7672 66 7700 2244
rect 7728 94 7756 2272
rect 7784 66 7812 2244
rect 7840 94 7868 2272
rect 7896 66 7924 2244
rect 7952 94 7980 2272
rect 8008 66 8036 2244
rect 8064 94 8092 2272
rect 8120 66 8148 2244
rect 8176 94 8204 2272
rect 8232 66 8260 2244
rect 8288 94 8316 2272
rect 8344 66 8372 2244
rect 8400 94 8428 2272
rect 8456 66 8484 2244
rect 8512 94 8540 2272
rect 8568 66 8596 2244
rect 8624 94 8652 2272
rect 8680 66 8708 2244
rect 8736 94 8764 2272
rect 8792 66 8820 2244
rect 8848 94 8876 2272
rect 8904 66 8932 2244
rect 8960 94 8988 2272
rect 9016 66 9044 2244
rect 9072 94 9100 2272
rect 9128 66 9156 2244
rect 9184 94 9212 2272
rect 9240 66 9268 2244
rect 9296 94 9324 2272
rect 9352 66 9380 2244
rect 9408 94 9436 2272
rect 9464 66 9492 2244
rect 9520 94 9548 2272
rect 9576 66 9604 2244
rect 9632 94 9660 2272
rect 9688 66 9716 2244
rect 9744 94 9772 2272
rect 9800 66 9828 2244
rect 9856 94 9884 2272
rect 9912 66 9940 2244
rect 9968 94 9996 2272
rect 10024 66 10052 2244
rect 10080 94 10108 2272
rect 10136 66 10164 2244
rect 10192 94 10220 2272
rect 10248 66 10276 2244
rect 10304 94 10332 2272
rect 10360 66 10388 2244
rect 10416 94 10444 2272
rect 10472 66 10500 2244
rect 10528 94 10556 2272
rect 10584 66 10612 2244
rect 10640 94 10668 2272
rect 10696 66 10724 2244
rect 10752 94 10780 2272
rect 10808 66 10836 2244
rect 10864 94 10892 2272
rect 10920 66 10948 2244
rect 10976 94 11004 2272
rect 11032 66 11060 2244
rect 11088 94 11146 2272
rect 0 59 11146 66
rect 0 7 24 59
rect 76 7 88 59
rect 140 50 236 59
rect 144 16 182 50
rect 216 16 236 50
rect 140 7 236 16
rect 288 7 300 59
rect 352 50 460 59
rect 360 16 398 50
rect 432 16 460 50
rect 352 7 460 16
rect 512 7 524 59
rect 576 50 684 59
rect 576 16 614 50
rect 648 16 684 50
rect 576 7 684 16
rect 736 7 748 59
rect 800 50 908 59
rect 800 16 830 50
rect 864 16 902 50
rect 800 7 908 16
rect 960 7 972 59
rect 1024 50 1132 59
rect 1184 50 1196 59
rect 1248 50 1356 59
rect 1408 50 1420 59
rect 1472 50 1580 59
rect 1632 50 1644 59
rect 1696 50 1804 59
rect 1856 50 1868 59
rect 1920 50 2028 59
rect 2080 50 2092 59
rect 2144 50 2252 59
rect 1024 16 1046 50
rect 1080 16 1118 50
rect 1184 16 1190 50
rect 1248 16 1262 50
rect 1296 16 1334 50
rect 1472 16 1478 50
rect 1512 16 1550 50
rect 1728 16 1766 50
rect 1800 16 1804 50
rect 1944 16 1982 50
rect 2016 16 2028 50
rect 2088 16 2092 50
rect 2160 16 2198 50
rect 2232 16 2252 50
rect 1024 7 1132 16
rect 1184 7 1196 16
rect 1248 7 1356 16
rect 1408 7 1420 16
rect 1472 7 1580 16
rect 1632 7 1644 16
rect 1696 7 1804 16
rect 1856 7 1868 16
rect 1920 7 2028 16
rect 2080 7 2092 16
rect 2144 7 2252 16
rect 2304 7 2316 59
rect 2368 50 2476 59
rect 2376 16 2414 50
rect 2448 16 2476 50
rect 2368 7 2476 16
rect 2528 7 2540 59
rect 2592 50 2700 59
rect 2592 16 2630 50
rect 2664 16 2700 50
rect 2592 7 2700 16
rect 2752 7 2764 59
rect 2816 50 2924 59
rect 2816 16 2846 50
rect 2880 16 2918 50
rect 2816 7 2924 16
rect 2976 7 2988 59
rect 3040 50 3148 59
rect 3200 50 3212 59
rect 3264 50 3372 59
rect 3424 50 3436 59
rect 3488 50 3596 59
rect 3648 50 3660 59
rect 3712 50 3820 59
rect 3872 50 3884 59
rect 3936 50 4044 59
rect 4096 50 4108 59
rect 4160 50 4268 59
rect 3040 16 3062 50
rect 3096 16 3134 50
rect 3200 16 3206 50
rect 3264 16 3278 50
rect 3312 16 3350 50
rect 3488 16 3494 50
rect 3528 16 3566 50
rect 3744 16 3782 50
rect 3816 16 3820 50
rect 3960 16 3998 50
rect 4032 16 4044 50
rect 4104 16 4108 50
rect 4176 16 4214 50
rect 4248 16 4268 50
rect 3040 7 3148 16
rect 3200 7 3212 16
rect 3264 7 3372 16
rect 3424 7 3436 16
rect 3488 7 3596 16
rect 3648 7 3660 16
rect 3712 7 3820 16
rect 3872 7 3884 16
rect 3936 7 4044 16
rect 4096 7 4108 16
rect 4160 7 4268 16
rect 4320 7 4332 59
rect 4384 50 4492 59
rect 4392 16 4430 50
rect 4464 16 4492 50
rect 4384 7 4492 16
rect 4544 7 4556 59
rect 4608 50 4716 59
rect 4608 16 4646 50
rect 4680 16 4716 50
rect 4608 7 4716 16
rect 4768 7 4780 59
rect 4832 50 4940 59
rect 4832 16 4862 50
rect 4896 16 4934 50
rect 4832 7 4940 16
rect 4992 7 5004 59
rect 5056 50 5164 59
rect 5216 50 5228 59
rect 5280 50 5388 59
rect 5440 50 5452 59
rect 5504 50 5612 59
rect 5664 50 5676 59
rect 5728 50 5836 59
rect 5888 50 5900 59
rect 5952 50 6060 59
rect 6112 50 6124 59
rect 6176 50 6284 59
rect 5056 16 5078 50
rect 5112 16 5150 50
rect 5216 16 5222 50
rect 5280 16 5294 50
rect 5328 16 5366 50
rect 5504 16 5510 50
rect 5544 16 5582 50
rect 5760 16 5798 50
rect 5832 16 5836 50
rect 5976 16 6014 50
rect 6048 16 6060 50
rect 6120 16 6124 50
rect 6192 16 6230 50
rect 6264 16 6284 50
rect 5056 7 5164 16
rect 5216 7 5228 16
rect 5280 7 5388 16
rect 5440 7 5452 16
rect 5504 7 5612 16
rect 5664 7 5676 16
rect 5728 7 5836 16
rect 5888 7 5900 16
rect 5952 7 6060 16
rect 6112 7 6124 16
rect 6176 7 6284 16
rect 6336 7 6348 59
rect 6400 50 6508 59
rect 6408 16 6446 50
rect 6480 16 6508 50
rect 6400 7 6508 16
rect 6560 7 6572 59
rect 6624 50 6732 59
rect 6624 16 6662 50
rect 6696 16 6732 50
rect 6624 7 6732 16
rect 6784 7 6796 59
rect 6848 50 6956 59
rect 6848 16 6878 50
rect 6912 16 6950 50
rect 6848 7 6956 16
rect 7008 7 7020 59
rect 7072 50 7180 59
rect 7232 50 7244 59
rect 7296 50 7404 59
rect 7456 50 7468 59
rect 7520 50 7628 59
rect 7680 50 7692 59
rect 7744 50 7852 59
rect 7904 50 7916 59
rect 7968 50 8076 59
rect 8128 50 8140 59
rect 8192 50 8300 59
rect 7072 16 7094 50
rect 7128 16 7166 50
rect 7232 16 7238 50
rect 7296 16 7310 50
rect 7344 16 7382 50
rect 7520 16 7526 50
rect 7560 16 7598 50
rect 7776 16 7814 50
rect 7848 16 7852 50
rect 7992 16 8030 50
rect 8064 16 8076 50
rect 8136 16 8140 50
rect 8208 16 8246 50
rect 8280 16 8300 50
rect 7072 7 7180 16
rect 7232 7 7244 16
rect 7296 7 7404 16
rect 7456 7 7468 16
rect 7520 7 7628 16
rect 7680 7 7692 16
rect 7744 7 7852 16
rect 7904 7 7916 16
rect 7968 7 8076 16
rect 8128 7 8140 16
rect 8192 7 8300 16
rect 8352 7 8364 59
rect 8416 50 8524 59
rect 8424 16 8462 50
rect 8496 16 8524 50
rect 8416 7 8524 16
rect 8576 7 8588 59
rect 8640 50 8748 59
rect 8640 16 8678 50
rect 8712 16 8748 50
rect 8640 7 8748 16
rect 8800 7 8812 59
rect 8864 50 8972 59
rect 8864 16 8894 50
rect 8928 16 8966 50
rect 8864 7 8972 16
rect 9024 7 9036 59
rect 9088 50 9196 59
rect 9248 50 9260 59
rect 9312 50 9420 59
rect 9472 50 9484 59
rect 9536 50 9644 59
rect 9696 50 9708 59
rect 9760 50 9868 59
rect 9920 50 9932 59
rect 9984 50 10092 59
rect 10144 50 10156 59
rect 10208 50 10316 59
rect 9088 16 9110 50
rect 9144 16 9182 50
rect 9248 16 9254 50
rect 9312 16 9326 50
rect 9360 16 9398 50
rect 9536 16 9542 50
rect 9576 16 9614 50
rect 9792 16 9830 50
rect 9864 16 9868 50
rect 10008 16 10046 50
rect 10080 16 10092 50
rect 10152 16 10156 50
rect 10224 16 10262 50
rect 10296 16 10316 50
rect 9088 7 9196 16
rect 9248 7 9260 16
rect 9312 7 9420 16
rect 9472 7 9484 16
rect 9536 7 9644 16
rect 9696 7 9708 16
rect 9760 7 9868 16
rect 9920 7 9932 16
rect 9984 7 10092 16
rect 10144 7 10156 16
rect 10208 7 10316 16
rect 10368 7 10380 59
rect 10432 50 10540 59
rect 10440 16 10478 50
rect 10512 16 10540 50
rect 10432 7 10540 16
rect 10592 7 10604 59
rect 10656 50 10764 59
rect 10656 16 10694 50
rect 10728 16 10764 50
rect 10656 7 10764 16
rect 10816 7 10828 59
rect 10880 50 10988 59
rect 10880 16 10910 50
rect 10944 16 10982 50
rect 10880 7 10988 16
rect 11040 7 11052 59
rect 11104 7 11146 59
rect 0 0 11146 7
<< via1 >>
rect 68 2322 120 2331
rect 132 2322 184 2331
rect 292 2322 344 2331
rect 356 2322 408 2331
rect 516 2322 568 2331
rect 580 2322 632 2331
rect 740 2322 792 2331
rect 68 2288 72 2322
rect 72 2288 110 2322
rect 110 2288 120 2322
rect 132 2288 144 2322
rect 144 2288 182 2322
rect 182 2288 184 2322
rect 292 2288 326 2322
rect 326 2288 344 2322
rect 356 2288 360 2322
rect 360 2288 398 2322
rect 398 2288 408 2322
rect 516 2288 542 2322
rect 542 2288 568 2322
rect 580 2288 614 2322
rect 614 2288 632 2322
rect 740 2288 758 2322
rect 758 2288 792 2322
rect 68 2279 120 2288
rect 132 2279 184 2288
rect 292 2279 344 2288
rect 356 2279 408 2288
rect 516 2279 568 2288
rect 580 2279 632 2288
rect 740 2279 792 2288
rect 804 2322 856 2331
rect 964 2322 1016 2331
rect 804 2288 830 2322
rect 830 2288 856 2322
rect 964 2288 974 2322
rect 974 2288 1008 2322
rect 1008 2288 1016 2322
rect 804 2279 856 2288
rect 964 2279 1016 2288
rect 1028 2322 1080 2331
rect 1188 2322 1240 2331
rect 1028 2288 1046 2322
rect 1046 2288 1080 2322
rect 1188 2288 1190 2322
rect 1190 2288 1224 2322
rect 1224 2288 1240 2322
rect 1028 2279 1080 2288
rect 1188 2279 1240 2288
rect 1252 2322 1304 2331
rect 1412 2322 1464 2331
rect 1252 2288 1262 2322
rect 1262 2288 1296 2322
rect 1296 2288 1304 2322
rect 1412 2288 1440 2322
rect 1440 2288 1464 2322
rect 1252 2279 1304 2288
rect 1412 2279 1464 2288
rect 1476 2322 1528 2331
rect 1636 2322 1688 2331
rect 1700 2322 1752 2331
rect 1860 2322 1912 2331
rect 1924 2322 1976 2331
rect 2084 2322 2136 2331
rect 2148 2322 2200 2331
rect 2308 2322 2360 2331
rect 2372 2322 2424 2331
rect 2532 2322 2584 2331
rect 2596 2322 2648 2331
rect 2756 2322 2808 2331
rect 1476 2288 1478 2322
rect 1478 2288 1512 2322
rect 1512 2288 1528 2322
rect 1636 2288 1656 2322
rect 1656 2288 1688 2322
rect 1700 2288 1728 2322
rect 1728 2288 1752 2322
rect 1860 2288 1872 2322
rect 1872 2288 1910 2322
rect 1910 2288 1912 2322
rect 1924 2288 1944 2322
rect 1944 2288 1976 2322
rect 2084 2288 2088 2322
rect 2088 2288 2126 2322
rect 2126 2288 2136 2322
rect 2148 2288 2160 2322
rect 2160 2288 2198 2322
rect 2198 2288 2200 2322
rect 2308 2288 2342 2322
rect 2342 2288 2360 2322
rect 2372 2288 2376 2322
rect 2376 2288 2414 2322
rect 2414 2288 2424 2322
rect 2532 2288 2558 2322
rect 2558 2288 2584 2322
rect 2596 2288 2630 2322
rect 2630 2288 2648 2322
rect 2756 2288 2774 2322
rect 2774 2288 2808 2322
rect 1476 2279 1528 2288
rect 1636 2279 1688 2288
rect 1700 2279 1752 2288
rect 1860 2279 1912 2288
rect 1924 2279 1976 2288
rect 2084 2279 2136 2288
rect 2148 2279 2200 2288
rect 2308 2279 2360 2288
rect 2372 2279 2424 2288
rect 2532 2279 2584 2288
rect 2596 2279 2648 2288
rect 2756 2279 2808 2288
rect 2820 2322 2872 2331
rect 2980 2322 3032 2331
rect 2820 2288 2846 2322
rect 2846 2288 2872 2322
rect 2980 2288 2990 2322
rect 2990 2288 3024 2322
rect 3024 2288 3032 2322
rect 2820 2279 2872 2288
rect 2980 2279 3032 2288
rect 3044 2322 3096 2331
rect 3204 2322 3256 2331
rect 3044 2288 3062 2322
rect 3062 2288 3096 2322
rect 3204 2288 3206 2322
rect 3206 2288 3240 2322
rect 3240 2288 3256 2322
rect 3044 2279 3096 2288
rect 3204 2279 3256 2288
rect 3268 2322 3320 2331
rect 3428 2322 3480 2331
rect 3268 2288 3278 2322
rect 3278 2288 3312 2322
rect 3312 2288 3320 2322
rect 3428 2288 3456 2322
rect 3456 2288 3480 2322
rect 3268 2279 3320 2288
rect 3428 2279 3480 2288
rect 3492 2322 3544 2331
rect 3652 2322 3704 2331
rect 3716 2322 3768 2331
rect 3876 2322 3928 2331
rect 3940 2322 3992 2331
rect 4100 2322 4152 2331
rect 4164 2322 4216 2331
rect 4324 2322 4376 2331
rect 4388 2322 4440 2331
rect 4548 2322 4600 2331
rect 4612 2322 4664 2331
rect 4772 2322 4824 2331
rect 3492 2288 3494 2322
rect 3494 2288 3528 2322
rect 3528 2288 3544 2322
rect 3652 2288 3672 2322
rect 3672 2288 3704 2322
rect 3716 2288 3744 2322
rect 3744 2288 3768 2322
rect 3876 2288 3888 2322
rect 3888 2288 3926 2322
rect 3926 2288 3928 2322
rect 3940 2288 3960 2322
rect 3960 2288 3992 2322
rect 4100 2288 4104 2322
rect 4104 2288 4142 2322
rect 4142 2288 4152 2322
rect 4164 2288 4176 2322
rect 4176 2288 4214 2322
rect 4214 2288 4216 2322
rect 4324 2288 4358 2322
rect 4358 2288 4376 2322
rect 4388 2288 4392 2322
rect 4392 2288 4430 2322
rect 4430 2288 4440 2322
rect 4548 2288 4574 2322
rect 4574 2288 4600 2322
rect 4612 2288 4646 2322
rect 4646 2288 4664 2322
rect 4772 2288 4790 2322
rect 4790 2288 4824 2322
rect 3492 2279 3544 2288
rect 3652 2279 3704 2288
rect 3716 2279 3768 2288
rect 3876 2279 3928 2288
rect 3940 2279 3992 2288
rect 4100 2279 4152 2288
rect 4164 2279 4216 2288
rect 4324 2279 4376 2288
rect 4388 2279 4440 2288
rect 4548 2279 4600 2288
rect 4612 2279 4664 2288
rect 4772 2279 4824 2288
rect 4836 2322 4888 2331
rect 4996 2322 5048 2331
rect 4836 2288 4862 2322
rect 4862 2288 4888 2322
rect 4996 2288 5006 2322
rect 5006 2288 5040 2322
rect 5040 2288 5048 2322
rect 4836 2279 4888 2288
rect 4996 2279 5048 2288
rect 5060 2322 5112 2331
rect 5220 2322 5272 2331
rect 5060 2288 5078 2322
rect 5078 2288 5112 2322
rect 5220 2288 5222 2322
rect 5222 2288 5256 2322
rect 5256 2288 5272 2322
rect 5060 2279 5112 2288
rect 5220 2279 5272 2288
rect 5284 2322 5336 2331
rect 5444 2322 5496 2331
rect 5284 2288 5294 2322
rect 5294 2288 5328 2322
rect 5328 2288 5336 2322
rect 5444 2288 5472 2322
rect 5472 2288 5496 2322
rect 5284 2279 5336 2288
rect 5444 2279 5496 2288
rect 5508 2322 5560 2331
rect 5668 2322 5720 2331
rect 5732 2322 5784 2331
rect 5892 2322 5944 2331
rect 5956 2322 6008 2331
rect 6116 2322 6168 2331
rect 6180 2322 6232 2331
rect 6340 2322 6392 2331
rect 6404 2322 6456 2331
rect 6564 2322 6616 2331
rect 6628 2322 6680 2331
rect 6788 2322 6840 2331
rect 5508 2288 5510 2322
rect 5510 2288 5544 2322
rect 5544 2288 5560 2322
rect 5668 2288 5688 2322
rect 5688 2288 5720 2322
rect 5732 2288 5760 2322
rect 5760 2288 5784 2322
rect 5892 2288 5904 2322
rect 5904 2288 5942 2322
rect 5942 2288 5944 2322
rect 5956 2288 5976 2322
rect 5976 2288 6008 2322
rect 6116 2288 6120 2322
rect 6120 2288 6158 2322
rect 6158 2288 6168 2322
rect 6180 2288 6192 2322
rect 6192 2288 6230 2322
rect 6230 2288 6232 2322
rect 6340 2288 6374 2322
rect 6374 2288 6392 2322
rect 6404 2288 6408 2322
rect 6408 2288 6446 2322
rect 6446 2288 6456 2322
rect 6564 2288 6590 2322
rect 6590 2288 6616 2322
rect 6628 2288 6662 2322
rect 6662 2288 6680 2322
rect 6788 2288 6806 2322
rect 6806 2288 6840 2322
rect 5508 2279 5560 2288
rect 5668 2279 5720 2288
rect 5732 2279 5784 2288
rect 5892 2279 5944 2288
rect 5956 2279 6008 2288
rect 6116 2279 6168 2288
rect 6180 2279 6232 2288
rect 6340 2279 6392 2288
rect 6404 2279 6456 2288
rect 6564 2279 6616 2288
rect 6628 2279 6680 2288
rect 6788 2279 6840 2288
rect 6852 2322 6904 2331
rect 7012 2322 7064 2331
rect 6852 2288 6878 2322
rect 6878 2288 6904 2322
rect 7012 2288 7022 2322
rect 7022 2288 7056 2322
rect 7056 2288 7064 2322
rect 6852 2279 6904 2288
rect 7012 2279 7064 2288
rect 7076 2322 7128 2331
rect 7236 2322 7288 2331
rect 7076 2288 7094 2322
rect 7094 2288 7128 2322
rect 7236 2288 7238 2322
rect 7238 2288 7272 2322
rect 7272 2288 7288 2322
rect 7076 2279 7128 2288
rect 7236 2279 7288 2288
rect 7300 2322 7352 2331
rect 7460 2322 7512 2331
rect 7300 2288 7310 2322
rect 7310 2288 7344 2322
rect 7344 2288 7352 2322
rect 7460 2288 7488 2322
rect 7488 2288 7512 2322
rect 7300 2279 7352 2288
rect 7460 2279 7512 2288
rect 7524 2322 7576 2331
rect 7684 2322 7736 2331
rect 7748 2322 7800 2331
rect 7908 2322 7960 2331
rect 7972 2322 8024 2331
rect 8132 2322 8184 2331
rect 8196 2322 8248 2331
rect 8356 2322 8408 2331
rect 8420 2322 8472 2331
rect 8580 2322 8632 2331
rect 8644 2322 8696 2331
rect 8804 2322 8856 2331
rect 7524 2288 7526 2322
rect 7526 2288 7560 2322
rect 7560 2288 7576 2322
rect 7684 2288 7704 2322
rect 7704 2288 7736 2322
rect 7748 2288 7776 2322
rect 7776 2288 7800 2322
rect 7908 2288 7920 2322
rect 7920 2288 7958 2322
rect 7958 2288 7960 2322
rect 7972 2288 7992 2322
rect 7992 2288 8024 2322
rect 8132 2288 8136 2322
rect 8136 2288 8174 2322
rect 8174 2288 8184 2322
rect 8196 2288 8208 2322
rect 8208 2288 8246 2322
rect 8246 2288 8248 2322
rect 8356 2288 8390 2322
rect 8390 2288 8408 2322
rect 8420 2288 8424 2322
rect 8424 2288 8462 2322
rect 8462 2288 8472 2322
rect 8580 2288 8606 2322
rect 8606 2288 8632 2322
rect 8644 2288 8678 2322
rect 8678 2288 8696 2322
rect 8804 2288 8822 2322
rect 8822 2288 8856 2322
rect 7524 2279 7576 2288
rect 7684 2279 7736 2288
rect 7748 2279 7800 2288
rect 7908 2279 7960 2288
rect 7972 2279 8024 2288
rect 8132 2279 8184 2288
rect 8196 2279 8248 2288
rect 8356 2279 8408 2288
rect 8420 2279 8472 2288
rect 8580 2279 8632 2288
rect 8644 2279 8696 2288
rect 8804 2279 8856 2288
rect 8868 2322 8920 2331
rect 9028 2322 9080 2331
rect 8868 2288 8894 2322
rect 8894 2288 8920 2322
rect 9028 2288 9038 2322
rect 9038 2288 9072 2322
rect 9072 2288 9080 2322
rect 8868 2279 8920 2288
rect 9028 2279 9080 2288
rect 9092 2322 9144 2331
rect 9252 2322 9304 2331
rect 9092 2288 9110 2322
rect 9110 2288 9144 2322
rect 9252 2288 9254 2322
rect 9254 2288 9288 2322
rect 9288 2288 9304 2322
rect 9092 2279 9144 2288
rect 9252 2279 9304 2288
rect 9316 2322 9368 2331
rect 9476 2322 9528 2331
rect 9316 2288 9326 2322
rect 9326 2288 9360 2322
rect 9360 2288 9368 2322
rect 9476 2288 9504 2322
rect 9504 2288 9528 2322
rect 9316 2279 9368 2288
rect 9476 2279 9528 2288
rect 9540 2322 9592 2331
rect 9700 2322 9752 2331
rect 9764 2322 9816 2331
rect 9924 2322 9976 2331
rect 9988 2322 10040 2331
rect 10148 2322 10200 2331
rect 10212 2322 10264 2331
rect 10372 2322 10424 2331
rect 10436 2322 10488 2331
rect 10596 2322 10648 2331
rect 10660 2322 10712 2331
rect 10820 2322 10872 2331
rect 9540 2288 9542 2322
rect 9542 2288 9576 2322
rect 9576 2288 9592 2322
rect 9700 2288 9720 2322
rect 9720 2288 9752 2322
rect 9764 2288 9792 2322
rect 9792 2288 9816 2322
rect 9924 2288 9936 2322
rect 9936 2288 9974 2322
rect 9974 2288 9976 2322
rect 9988 2288 10008 2322
rect 10008 2288 10040 2322
rect 10148 2288 10152 2322
rect 10152 2288 10190 2322
rect 10190 2288 10200 2322
rect 10212 2288 10224 2322
rect 10224 2288 10262 2322
rect 10262 2288 10264 2322
rect 10372 2288 10406 2322
rect 10406 2288 10424 2322
rect 10436 2288 10440 2322
rect 10440 2288 10478 2322
rect 10478 2288 10488 2322
rect 10596 2288 10622 2322
rect 10622 2288 10648 2322
rect 10660 2288 10694 2322
rect 10694 2288 10712 2322
rect 10820 2288 10838 2322
rect 10838 2288 10872 2322
rect 9540 2279 9592 2288
rect 9700 2279 9752 2288
rect 9764 2279 9816 2288
rect 9924 2279 9976 2288
rect 9988 2279 10040 2288
rect 10148 2279 10200 2288
rect 10212 2279 10264 2288
rect 10372 2279 10424 2288
rect 10436 2279 10488 2288
rect 10596 2279 10648 2288
rect 10660 2279 10712 2288
rect 10820 2279 10872 2288
rect 10884 2322 10936 2331
rect 10884 2288 10910 2322
rect 10910 2288 10936 2322
rect 10884 2279 10936 2288
rect 24 50 76 59
rect 24 16 38 50
rect 38 16 72 50
rect 72 16 76 50
rect 24 7 76 16
rect 88 50 140 59
rect 236 50 288 59
rect 88 16 110 50
rect 110 16 140 50
rect 236 16 254 50
rect 254 16 288 50
rect 88 7 140 16
rect 236 7 288 16
rect 300 50 352 59
rect 460 50 512 59
rect 300 16 326 50
rect 326 16 352 50
rect 460 16 470 50
rect 470 16 504 50
rect 504 16 512 50
rect 300 7 352 16
rect 460 7 512 16
rect 524 50 576 59
rect 684 50 736 59
rect 524 16 542 50
rect 542 16 576 50
rect 684 16 686 50
rect 686 16 720 50
rect 720 16 736 50
rect 524 7 576 16
rect 684 7 736 16
rect 748 50 800 59
rect 908 50 960 59
rect 748 16 758 50
rect 758 16 792 50
rect 792 16 800 50
rect 908 16 936 50
rect 936 16 960 50
rect 748 7 800 16
rect 908 7 960 16
rect 972 50 1024 59
rect 1132 50 1184 59
rect 1196 50 1248 59
rect 1356 50 1408 59
rect 1420 50 1472 59
rect 1580 50 1632 59
rect 1644 50 1696 59
rect 1804 50 1856 59
rect 1868 50 1920 59
rect 2028 50 2080 59
rect 2092 50 2144 59
rect 2252 50 2304 59
rect 972 16 974 50
rect 974 16 1008 50
rect 1008 16 1024 50
rect 1132 16 1152 50
rect 1152 16 1184 50
rect 1196 16 1224 50
rect 1224 16 1248 50
rect 1356 16 1368 50
rect 1368 16 1406 50
rect 1406 16 1408 50
rect 1420 16 1440 50
rect 1440 16 1472 50
rect 1580 16 1584 50
rect 1584 16 1622 50
rect 1622 16 1632 50
rect 1644 16 1656 50
rect 1656 16 1694 50
rect 1694 16 1696 50
rect 1804 16 1838 50
rect 1838 16 1856 50
rect 1868 16 1872 50
rect 1872 16 1910 50
rect 1910 16 1920 50
rect 2028 16 2054 50
rect 2054 16 2080 50
rect 2092 16 2126 50
rect 2126 16 2144 50
rect 2252 16 2270 50
rect 2270 16 2304 50
rect 972 7 1024 16
rect 1132 7 1184 16
rect 1196 7 1248 16
rect 1356 7 1408 16
rect 1420 7 1472 16
rect 1580 7 1632 16
rect 1644 7 1696 16
rect 1804 7 1856 16
rect 1868 7 1920 16
rect 2028 7 2080 16
rect 2092 7 2144 16
rect 2252 7 2304 16
rect 2316 50 2368 59
rect 2476 50 2528 59
rect 2316 16 2342 50
rect 2342 16 2368 50
rect 2476 16 2486 50
rect 2486 16 2520 50
rect 2520 16 2528 50
rect 2316 7 2368 16
rect 2476 7 2528 16
rect 2540 50 2592 59
rect 2700 50 2752 59
rect 2540 16 2558 50
rect 2558 16 2592 50
rect 2700 16 2702 50
rect 2702 16 2736 50
rect 2736 16 2752 50
rect 2540 7 2592 16
rect 2700 7 2752 16
rect 2764 50 2816 59
rect 2924 50 2976 59
rect 2764 16 2774 50
rect 2774 16 2808 50
rect 2808 16 2816 50
rect 2924 16 2952 50
rect 2952 16 2976 50
rect 2764 7 2816 16
rect 2924 7 2976 16
rect 2988 50 3040 59
rect 3148 50 3200 59
rect 3212 50 3264 59
rect 3372 50 3424 59
rect 3436 50 3488 59
rect 3596 50 3648 59
rect 3660 50 3712 59
rect 3820 50 3872 59
rect 3884 50 3936 59
rect 4044 50 4096 59
rect 4108 50 4160 59
rect 4268 50 4320 59
rect 2988 16 2990 50
rect 2990 16 3024 50
rect 3024 16 3040 50
rect 3148 16 3168 50
rect 3168 16 3200 50
rect 3212 16 3240 50
rect 3240 16 3264 50
rect 3372 16 3384 50
rect 3384 16 3422 50
rect 3422 16 3424 50
rect 3436 16 3456 50
rect 3456 16 3488 50
rect 3596 16 3600 50
rect 3600 16 3638 50
rect 3638 16 3648 50
rect 3660 16 3672 50
rect 3672 16 3710 50
rect 3710 16 3712 50
rect 3820 16 3854 50
rect 3854 16 3872 50
rect 3884 16 3888 50
rect 3888 16 3926 50
rect 3926 16 3936 50
rect 4044 16 4070 50
rect 4070 16 4096 50
rect 4108 16 4142 50
rect 4142 16 4160 50
rect 4268 16 4286 50
rect 4286 16 4320 50
rect 2988 7 3040 16
rect 3148 7 3200 16
rect 3212 7 3264 16
rect 3372 7 3424 16
rect 3436 7 3488 16
rect 3596 7 3648 16
rect 3660 7 3712 16
rect 3820 7 3872 16
rect 3884 7 3936 16
rect 4044 7 4096 16
rect 4108 7 4160 16
rect 4268 7 4320 16
rect 4332 50 4384 59
rect 4492 50 4544 59
rect 4332 16 4358 50
rect 4358 16 4384 50
rect 4492 16 4502 50
rect 4502 16 4536 50
rect 4536 16 4544 50
rect 4332 7 4384 16
rect 4492 7 4544 16
rect 4556 50 4608 59
rect 4716 50 4768 59
rect 4556 16 4574 50
rect 4574 16 4608 50
rect 4716 16 4718 50
rect 4718 16 4752 50
rect 4752 16 4768 50
rect 4556 7 4608 16
rect 4716 7 4768 16
rect 4780 50 4832 59
rect 4940 50 4992 59
rect 4780 16 4790 50
rect 4790 16 4824 50
rect 4824 16 4832 50
rect 4940 16 4968 50
rect 4968 16 4992 50
rect 4780 7 4832 16
rect 4940 7 4992 16
rect 5004 50 5056 59
rect 5164 50 5216 59
rect 5228 50 5280 59
rect 5388 50 5440 59
rect 5452 50 5504 59
rect 5612 50 5664 59
rect 5676 50 5728 59
rect 5836 50 5888 59
rect 5900 50 5952 59
rect 6060 50 6112 59
rect 6124 50 6176 59
rect 6284 50 6336 59
rect 5004 16 5006 50
rect 5006 16 5040 50
rect 5040 16 5056 50
rect 5164 16 5184 50
rect 5184 16 5216 50
rect 5228 16 5256 50
rect 5256 16 5280 50
rect 5388 16 5400 50
rect 5400 16 5438 50
rect 5438 16 5440 50
rect 5452 16 5472 50
rect 5472 16 5504 50
rect 5612 16 5616 50
rect 5616 16 5654 50
rect 5654 16 5664 50
rect 5676 16 5688 50
rect 5688 16 5726 50
rect 5726 16 5728 50
rect 5836 16 5870 50
rect 5870 16 5888 50
rect 5900 16 5904 50
rect 5904 16 5942 50
rect 5942 16 5952 50
rect 6060 16 6086 50
rect 6086 16 6112 50
rect 6124 16 6158 50
rect 6158 16 6176 50
rect 6284 16 6302 50
rect 6302 16 6336 50
rect 5004 7 5056 16
rect 5164 7 5216 16
rect 5228 7 5280 16
rect 5388 7 5440 16
rect 5452 7 5504 16
rect 5612 7 5664 16
rect 5676 7 5728 16
rect 5836 7 5888 16
rect 5900 7 5952 16
rect 6060 7 6112 16
rect 6124 7 6176 16
rect 6284 7 6336 16
rect 6348 50 6400 59
rect 6508 50 6560 59
rect 6348 16 6374 50
rect 6374 16 6400 50
rect 6508 16 6518 50
rect 6518 16 6552 50
rect 6552 16 6560 50
rect 6348 7 6400 16
rect 6508 7 6560 16
rect 6572 50 6624 59
rect 6732 50 6784 59
rect 6572 16 6590 50
rect 6590 16 6624 50
rect 6732 16 6734 50
rect 6734 16 6768 50
rect 6768 16 6784 50
rect 6572 7 6624 16
rect 6732 7 6784 16
rect 6796 50 6848 59
rect 6956 50 7008 59
rect 6796 16 6806 50
rect 6806 16 6840 50
rect 6840 16 6848 50
rect 6956 16 6984 50
rect 6984 16 7008 50
rect 6796 7 6848 16
rect 6956 7 7008 16
rect 7020 50 7072 59
rect 7180 50 7232 59
rect 7244 50 7296 59
rect 7404 50 7456 59
rect 7468 50 7520 59
rect 7628 50 7680 59
rect 7692 50 7744 59
rect 7852 50 7904 59
rect 7916 50 7968 59
rect 8076 50 8128 59
rect 8140 50 8192 59
rect 8300 50 8352 59
rect 7020 16 7022 50
rect 7022 16 7056 50
rect 7056 16 7072 50
rect 7180 16 7200 50
rect 7200 16 7232 50
rect 7244 16 7272 50
rect 7272 16 7296 50
rect 7404 16 7416 50
rect 7416 16 7454 50
rect 7454 16 7456 50
rect 7468 16 7488 50
rect 7488 16 7520 50
rect 7628 16 7632 50
rect 7632 16 7670 50
rect 7670 16 7680 50
rect 7692 16 7704 50
rect 7704 16 7742 50
rect 7742 16 7744 50
rect 7852 16 7886 50
rect 7886 16 7904 50
rect 7916 16 7920 50
rect 7920 16 7958 50
rect 7958 16 7968 50
rect 8076 16 8102 50
rect 8102 16 8128 50
rect 8140 16 8174 50
rect 8174 16 8192 50
rect 8300 16 8318 50
rect 8318 16 8352 50
rect 7020 7 7072 16
rect 7180 7 7232 16
rect 7244 7 7296 16
rect 7404 7 7456 16
rect 7468 7 7520 16
rect 7628 7 7680 16
rect 7692 7 7744 16
rect 7852 7 7904 16
rect 7916 7 7968 16
rect 8076 7 8128 16
rect 8140 7 8192 16
rect 8300 7 8352 16
rect 8364 50 8416 59
rect 8524 50 8576 59
rect 8364 16 8390 50
rect 8390 16 8416 50
rect 8524 16 8534 50
rect 8534 16 8568 50
rect 8568 16 8576 50
rect 8364 7 8416 16
rect 8524 7 8576 16
rect 8588 50 8640 59
rect 8748 50 8800 59
rect 8588 16 8606 50
rect 8606 16 8640 50
rect 8748 16 8750 50
rect 8750 16 8784 50
rect 8784 16 8800 50
rect 8588 7 8640 16
rect 8748 7 8800 16
rect 8812 50 8864 59
rect 8972 50 9024 59
rect 8812 16 8822 50
rect 8822 16 8856 50
rect 8856 16 8864 50
rect 8972 16 9000 50
rect 9000 16 9024 50
rect 8812 7 8864 16
rect 8972 7 9024 16
rect 9036 50 9088 59
rect 9196 50 9248 59
rect 9260 50 9312 59
rect 9420 50 9472 59
rect 9484 50 9536 59
rect 9644 50 9696 59
rect 9708 50 9760 59
rect 9868 50 9920 59
rect 9932 50 9984 59
rect 10092 50 10144 59
rect 10156 50 10208 59
rect 10316 50 10368 59
rect 9036 16 9038 50
rect 9038 16 9072 50
rect 9072 16 9088 50
rect 9196 16 9216 50
rect 9216 16 9248 50
rect 9260 16 9288 50
rect 9288 16 9312 50
rect 9420 16 9432 50
rect 9432 16 9470 50
rect 9470 16 9472 50
rect 9484 16 9504 50
rect 9504 16 9536 50
rect 9644 16 9648 50
rect 9648 16 9686 50
rect 9686 16 9696 50
rect 9708 16 9720 50
rect 9720 16 9758 50
rect 9758 16 9760 50
rect 9868 16 9902 50
rect 9902 16 9920 50
rect 9932 16 9936 50
rect 9936 16 9974 50
rect 9974 16 9984 50
rect 10092 16 10118 50
rect 10118 16 10144 50
rect 10156 16 10190 50
rect 10190 16 10208 50
rect 10316 16 10334 50
rect 10334 16 10368 50
rect 9036 7 9088 16
rect 9196 7 9248 16
rect 9260 7 9312 16
rect 9420 7 9472 16
rect 9484 7 9536 16
rect 9644 7 9696 16
rect 9708 7 9760 16
rect 9868 7 9920 16
rect 9932 7 9984 16
rect 10092 7 10144 16
rect 10156 7 10208 16
rect 10316 7 10368 16
rect 10380 50 10432 59
rect 10540 50 10592 59
rect 10380 16 10406 50
rect 10406 16 10432 50
rect 10540 16 10550 50
rect 10550 16 10584 50
rect 10584 16 10592 50
rect 10380 7 10432 16
rect 10540 7 10592 16
rect 10604 50 10656 59
rect 10764 50 10816 59
rect 10604 16 10622 50
rect 10622 16 10656 50
rect 10764 16 10766 50
rect 10766 16 10800 50
rect 10800 16 10816 50
rect 10604 7 10656 16
rect 10764 7 10816 16
rect 10828 50 10880 59
rect 10988 50 11040 59
rect 10828 16 10838 50
rect 10838 16 10872 50
rect 10872 16 10880 50
rect 10988 16 11016 50
rect 11016 16 11040 50
rect 10828 7 10880 16
rect 10988 7 11040 16
rect 11052 50 11104 59
rect 11052 16 11054 50
rect 11054 16 11088 50
rect 11088 16 11104 50
rect 11052 7 11104 16
<< metal2 >>
rect 0 66 28 2338
rect 56 2333 196 2338
rect 56 2331 98 2333
rect 154 2331 196 2333
rect 56 2279 68 2331
rect 184 2279 196 2331
rect 56 2277 98 2279
rect 154 2277 196 2279
rect 56 2272 196 2277
rect 56 94 84 2272
rect 112 66 140 2244
rect 0 61 140 66
rect 0 59 42 61
rect 98 59 140 61
rect 0 7 24 59
rect 0 5 42 7
rect 98 5 140 7
rect 0 0 140 5
rect 168 0 196 2272
rect 224 66 252 2338
rect 280 2333 420 2338
rect 280 2331 322 2333
rect 378 2331 420 2333
rect 280 2279 292 2331
rect 408 2279 420 2331
rect 280 2277 322 2279
rect 378 2277 420 2279
rect 280 2272 420 2277
rect 280 94 308 2272
rect 336 66 364 2244
rect 224 61 364 66
rect 224 59 266 61
rect 322 59 364 61
rect 224 7 236 59
rect 352 7 364 59
rect 224 5 266 7
rect 322 5 364 7
rect 224 0 364 5
rect 392 0 420 2272
rect 448 66 476 2338
rect 504 2333 644 2338
rect 504 2331 546 2333
rect 602 2331 644 2333
rect 504 2279 516 2331
rect 632 2279 644 2331
rect 504 2277 546 2279
rect 602 2277 644 2279
rect 504 2272 644 2277
rect 504 94 532 2272
rect 560 66 588 2244
rect 448 61 588 66
rect 448 59 490 61
rect 546 59 588 61
rect 448 7 460 59
rect 576 7 588 59
rect 448 5 490 7
rect 546 5 588 7
rect 448 0 588 5
rect 616 0 644 2272
rect 672 66 700 2338
rect 728 2333 868 2338
rect 728 2331 770 2333
rect 826 2331 868 2333
rect 728 2279 740 2331
rect 856 2279 868 2331
rect 728 2277 770 2279
rect 826 2277 868 2279
rect 728 2272 868 2277
rect 728 94 756 2272
rect 784 66 812 2244
rect 672 61 812 66
rect 672 59 714 61
rect 770 59 812 61
rect 672 7 684 59
rect 800 7 812 59
rect 672 5 714 7
rect 770 5 812 7
rect 672 0 812 5
rect 840 0 868 2272
rect 896 66 924 2338
rect 952 2333 1092 2338
rect 952 2331 994 2333
rect 1050 2331 1092 2333
rect 952 2279 964 2331
rect 1080 2279 1092 2331
rect 952 2277 994 2279
rect 1050 2277 1092 2279
rect 952 2272 1092 2277
rect 952 94 980 2272
rect 1008 66 1036 2244
rect 896 61 1036 66
rect 896 59 938 61
rect 994 59 1036 61
rect 896 7 908 59
rect 1024 7 1036 59
rect 896 5 938 7
rect 994 5 1036 7
rect 896 0 1036 5
rect 1064 0 1092 2272
rect 1120 66 1148 2338
rect 1176 2333 1316 2338
rect 1176 2331 1218 2333
rect 1274 2331 1316 2333
rect 1176 2279 1188 2331
rect 1304 2279 1316 2331
rect 1176 2277 1218 2279
rect 1274 2277 1316 2279
rect 1176 2272 1316 2277
rect 1176 94 1204 2272
rect 1232 66 1260 2244
rect 1120 61 1260 66
rect 1120 59 1162 61
rect 1218 59 1260 61
rect 1120 7 1132 59
rect 1248 7 1260 59
rect 1120 5 1162 7
rect 1218 5 1260 7
rect 1120 0 1260 5
rect 1288 0 1316 2272
rect 1344 66 1372 2338
rect 1400 2333 1540 2338
rect 1400 2331 1442 2333
rect 1498 2331 1540 2333
rect 1400 2279 1412 2331
rect 1528 2279 1540 2331
rect 1400 2277 1442 2279
rect 1498 2277 1540 2279
rect 1400 2272 1540 2277
rect 1400 94 1428 2272
rect 1456 66 1484 2244
rect 1344 61 1484 66
rect 1344 59 1386 61
rect 1442 59 1484 61
rect 1344 7 1356 59
rect 1472 7 1484 59
rect 1344 5 1386 7
rect 1442 5 1484 7
rect 1344 0 1484 5
rect 1512 0 1540 2272
rect 1568 66 1596 2338
rect 1624 2333 1764 2338
rect 1624 2331 1666 2333
rect 1722 2331 1764 2333
rect 1624 2279 1636 2331
rect 1752 2279 1764 2331
rect 1624 2277 1666 2279
rect 1722 2277 1764 2279
rect 1624 2272 1764 2277
rect 1624 94 1652 2272
rect 1680 66 1708 2244
rect 1568 61 1708 66
rect 1568 59 1610 61
rect 1666 59 1708 61
rect 1568 7 1580 59
rect 1696 7 1708 59
rect 1568 5 1610 7
rect 1666 5 1708 7
rect 1568 0 1708 5
rect 1736 0 1764 2272
rect 1792 66 1820 2338
rect 1848 2333 1988 2338
rect 1848 2331 1890 2333
rect 1946 2331 1988 2333
rect 1848 2279 1860 2331
rect 1976 2279 1988 2331
rect 1848 2277 1890 2279
rect 1946 2277 1988 2279
rect 1848 2272 1988 2277
rect 1848 94 1876 2272
rect 1904 66 1932 2244
rect 1792 61 1932 66
rect 1792 59 1834 61
rect 1890 59 1932 61
rect 1792 7 1804 59
rect 1920 7 1932 59
rect 1792 5 1834 7
rect 1890 5 1932 7
rect 1792 0 1932 5
rect 1960 0 1988 2272
rect 2016 66 2044 2338
rect 2072 2333 2212 2338
rect 2072 2331 2114 2333
rect 2170 2331 2212 2333
rect 2072 2279 2084 2331
rect 2200 2279 2212 2331
rect 2072 2277 2114 2279
rect 2170 2277 2212 2279
rect 2072 2272 2212 2277
rect 2072 94 2100 2272
rect 2128 66 2156 2244
rect 2016 61 2156 66
rect 2016 59 2058 61
rect 2114 59 2156 61
rect 2016 7 2028 59
rect 2144 7 2156 59
rect 2016 5 2058 7
rect 2114 5 2156 7
rect 2016 0 2156 5
rect 2184 0 2212 2272
rect 2240 66 2268 2338
rect 2296 2333 2436 2338
rect 2296 2331 2338 2333
rect 2394 2331 2436 2333
rect 2296 2279 2308 2331
rect 2424 2279 2436 2331
rect 2296 2277 2338 2279
rect 2394 2277 2436 2279
rect 2296 2272 2436 2277
rect 2296 94 2324 2272
rect 2352 66 2380 2244
rect 2240 61 2380 66
rect 2240 59 2282 61
rect 2338 59 2380 61
rect 2240 7 2252 59
rect 2368 7 2380 59
rect 2240 5 2282 7
rect 2338 5 2380 7
rect 2240 0 2380 5
rect 2408 0 2436 2272
rect 2464 66 2492 2338
rect 2520 2333 2660 2338
rect 2520 2331 2562 2333
rect 2618 2331 2660 2333
rect 2520 2279 2532 2331
rect 2648 2279 2660 2331
rect 2520 2277 2562 2279
rect 2618 2277 2660 2279
rect 2520 2272 2660 2277
rect 2520 94 2548 2272
rect 2576 66 2604 2244
rect 2464 61 2604 66
rect 2464 59 2506 61
rect 2562 59 2604 61
rect 2464 7 2476 59
rect 2592 7 2604 59
rect 2464 5 2506 7
rect 2562 5 2604 7
rect 2464 0 2604 5
rect 2632 0 2660 2272
rect 2688 66 2716 2338
rect 2744 2333 2884 2338
rect 2744 2331 2786 2333
rect 2842 2331 2884 2333
rect 2744 2279 2756 2331
rect 2872 2279 2884 2331
rect 2744 2277 2786 2279
rect 2842 2277 2884 2279
rect 2744 2272 2884 2277
rect 2744 94 2772 2272
rect 2800 66 2828 2244
rect 2688 61 2828 66
rect 2688 59 2730 61
rect 2786 59 2828 61
rect 2688 7 2700 59
rect 2816 7 2828 59
rect 2688 5 2730 7
rect 2786 5 2828 7
rect 2688 0 2828 5
rect 2856 0 2884 2272
rect 2912 66 2940 2338
rect 2968 2333 3108 2338
rect 2968 2331 3010 2333
rect 3066 2331 3108 2333
rect 2968 2279 2980 2331
rect 3096 2279 3108 2331
rect 2968 2277 3010 2279
rect 3066 2277 3108 2279
rect 2968 2272 3108 2277
rect 2968 94 2996 2272
rect 3024 66 3052 2244
rect 2912 61 3052 66
rect 2912 59 2954 61
rect 3010 59 3052 61
rect 2912 7 2924 59
rect 3040 7 3052 59
rect 2912 5 2954 7
rect 3010 5 3052 7
rect 2912 0 3052 5
rect 3080 0 3108 2272
rect 3136 66 3164 2338
rect 3192 2333 3332 2338
rect 3192 2331 3234 2333
rect 3290 2331 3332 2333
rect 3192 2279 3204 2331
rect 3320 2279 3332 2331
rect 3192 2277 3234 2279
rect 3290 2277 3332 2279
rect 3192 2272 3332 2277
rect 3192 94 3220 2272
rect 3248 66 3276 2244
rect 3136 61 3276 66
rect 3136 59 3178 61
rect 3234 59 3276 61
rect 3136 7 3148 59
rect 3264 7 3276 59
rect 3136 5 3178 7
rect 3234 5 3276 7
rect 3136 0 3276 5
rect 3304 0 3332 2272
rect 3360 66 3388 2338
rect 3416 2333 3556 2338
rect 3416 2331 3458 2333
rect 3514 2331 3556 2333
rect 3416 2279 3428 2331
rect 3544 2279 3556 2331
rect 3416 2277 3458 2279
rect 3514 2277 3556 2279
rect 3416 2272 3556 2277
rect 3416 94 3444 2272
rect 3472 66 3500 2244
rect 3360 61 3500 66
rect 3360 59 3402 61
rect 3458 59 3500 61
rect 3360 7 3372 59
rect 3488 7 3500 59
rect 3360 5 3402 7
rect 3458 5 3500 7
rect 3360 0 3500 5
rect 3528 0 3556 2272
rect 3584 66 3612 2338
rect 3640 2333 3780 2338
rect 3640 2331 3682 2333
rect 3738 2331 3780 2333
rect 3640 2279 3652 2331
rect 3768 2279 3780 2331
rect 3640 2277 3682 2279
rect 3738 2277 3780 2279
rect 3640 2272 3780 2277
rect 3640 94 3668 2272
rect 3696 66 3724 2244
rect 3584 61 3724 66
rect 3584 59 3626 61
rect 3682 59 3724 61
rect 3584 7 3596 59
rect 3712 7 3724 59
rect 3584 5 3626 7
rect 3682 5 3724 7
rect 3584 0 3724 5
rect 3752 0 3780 2272
rect 3808 66 3836 2338
rect 3864 2333 4004 2338
rect 3864 2331 3906 2333
rect 3962 2331 4004 2333
rect 3864 2279 3876 2331
rect 3992 2279 4004 2331
rect 3864 2277 3906 2279
rect 3962 2277 4004 2279
rect 3864 2272 4004 2277
rect 3864 94 3892 2272
rect 3920 66 3948 2244
rect 3808 61 3948 66
rect 3808 59 3850 61
rect 3906 59 3948 61
rect 3808 7 3820 59
rect 3936 7 3948 59
rect 3808 5 3850 7
rect 3906 5 3948 7
rect 3808 0 3948 5
rect 3976 0 4004 2272
rect 4032 66 4060 2338
rect 4088 2333 4228 2338
rect 4088 2331 4130 2333
rect 4186 2331 4228 2333
rect 4088 2279 4100 2331
rect 4216 2279 4228 2331
rect 4088 2277 4130 2279
rect 4186 2277 4228 2279
rect 4088 2272 4228 2277
rect 4088 94 4116 2272
rect 4144 66 4172 2244
rect 4032 61 4172 66
rect 4032 59 4074 61
rect 4130 59 4172 61
rect 4032 7 4044 59
rect 4160 7 4172 59
rect 4032 5 4074 7
rect 4130 5 4172 7
rect 4032 0 4172 5
rect 4200 0 4228 2272
rect 4256 66 4284 2338
rect 4312 2333 4452 2338
rect 4312 2331 4354 2333
rect 4410 2331 4452 2333
rect 4312 2279 4324 2331
rect 4440 2279 4452 2331
rect 4312 2277 4354 2279
rect 4410 2277 4452 2279
rect 4312 2272 4452 2277
rect 4312 94 4340 2272
rect 4368 66 4396 2244
rect 4256 61 4396 66
rect 4256 59 4298 61
rect 4354 59 4396 61
rect 4256 7 4268 59
rect 4384 7 4396 59
rect 4256 5 4298 7
rect 4354 5 4396 7
rect 4256 0 4396 5
rect 4424 0 4452 2272
rect 4480 66 4508 2338
rect 4536 2333 4676 2338
rect 4536 2331 4578 2333
rect 4634 2331 4676 2333
rect 4536 2279 4548 2331
rect 4664 2279 4676 2331
rect 4536 2277 4578 2279
rect 4634 2277 4676 2279
rect 4536 2272 4676 2277
rect 4536 94 4564 2272
rect 4592 66 4620 2244
rect 4480 61 4620 66
rect 4480 59 4522 61
rect 4578 59 4620 61
rect 4480 7 4492 59
rect 4608 7 4620 59
rect 4480 5 4522 7
rect 4578 5 4620 7
rect 4480 0 4620 5
rect 4648 0 4676 2272
rect 4704 66 4732 2338
rect 4760 2333 4900 2338
rect 4760 2331 4802 2333
rect 4858 2331 4900 2333
rect 4760 2279 4772 2331
rect 4888 2279 4900 2331
rect 4760 2277 4802 2279
rect 4858 2277 4900 2279
rect 4760 2272 4900 2277
rect 4760 94 4788 2272
rect 4816 66 4844 2244
rect 4704 61 4844 66
rect 4704 59 4746 61
rect 4802 59 4844 61
rect 4704 7 4716 59
rect 4832 7 4844 59
rect 4704 5 4746 7
rect 4802 5 4844 7
rect 4704 0 4844 5
rect 4872 0 4900 2272
rect 4928 66 4956 2338
rect 4984 2333 5124 2338
rect 4984 2331 5026 2333
rect 5082 2331 5124 2333
rect 4984 2279 4996 2331
rect 5112 2279 5124 2331
rect 4984 2277 5026 2279
rect 5082 2277 5124 2279
rect 4984 2272 5124 2277
rect 4984 94 5012 2272
rect 5040 66 5068 2244
rect 4928 61 5068 66
rect 4928 59 4970 61
rect 5026 59 5068 61
rect 4928 7 4940 59
rect 5056 7 5068 59
rect 4928 5 4970 7
rect 5026 5 5068 7
rect 4928 0 5068 5
rect 5096 0 5124 2272
rect 5152 66 5180 2338
rect 5208 2333 5348 2338
rect 5208 2331 5250 2333
rect 5306 2331 5348 2333
rect 5208 2279 5220 2331
rect 5336 2279 5348 2331
rect 5208 2277 5250 2279
rect 5306 2277 5348 2279
rect 5208 2272 5348 2277
rect 5208 94 5236 2272
rect 5264 66 5292 2244
rect 5152 61 5292 66
rect 5152 59 5194 61
rect 5250 59 5292 61
rect 5152 7 5164 59
rect 5280 7 5292 59
rect 5152 5 5194 7
rect 5250 5 5292 7
rect 5152 0 5292 5
rect 5320 0 5348 2272
rect 5376 66 5404 2338
rect 5432 2333 5572 2338
rect 5432 2331 5474 2333
rect 5530 2331 5572 2333
rect 5432 2279 5444 2331
rect 5560 2279 5572 2331
rect 5432 2277 5474 2279
rect 5530 2277 5572 2279
rect 5432 2272 5572 2277
rect 5432 94 5460 2272
rect 5488 66 5516 2244
rect 5376 61 5516 66
rect 5376 59 5418 61
rect 5474 59 5516 61
rect 5376 7 5388 59
rect 5504 7 5516 59
rect 5376 5 5418 7
rect 5474 5 5516 7
rect 5376 0 5516 5
rect 5544 0 5572 2272
rect 5600 66 5628 2338
rect 5656 2333 5796 2338
rect 5656 2331 5698 2333
rect 5754 2331 5796 2333
rect 5656 2279 5668 2331
rect 5784 2279 5796 2331
rect 5656 2277 5698 2279
rect 5754 2277 5796 2279
rect 5656 2272 5796 2277
rect 5656 94 5684 2272
rect 5712 66 5740 2244
rect 5600 61 5740 66
rect 5600 59 5642 61
rect 5698 59 5740 61
rect 5600 7 5612 59
rect 5728 7 5740 59
rect 5600 5 5642 7
rect 5698 5 5740 7
rect 5600 0 5740 5
rect 5768 0 5796 2272
rect 5824 66 5852 2338
rect 5880 2333 6020 2338
rect 5880 2331 5922 2333
rect 5978 2331 6020 2333
rect 5880 2279 5892 2331
rect 6008 2279 6020 2331
rect 5880 2277 5922 2279
rect 5978 2277 6020 2279
rect 5880 2272 6020 2277
rect 5880 94 5908 2272
rect 5936 66 5964 2244
rect 5824 61 5964 66
rect 5824 59 5866 61
rect 5922 59 5964 61
rect 5824 7 5836 59
rect 5952 7 5964 59
rect 5824 5 5866 7
rect 5922 5 5964 7
rect 5824 0 5964 5
rect 5992 0 6020 2272
rect 6048 66 6076 2338
rect 6104 2333 6244 2338
rect 6104 2331 6146 2333
rect 6202 2331 6244 2333
rect 6104 2279 6116 2331
rect 6232 2279 6244 2331
rect 6104 2277 6146 2279
rect 6202 2277 6244 2279
rect 6104 2272 6244 2277
rect 6104 94 6132 2272
rect 6160 66 6188 2244
rect 6048 61 6188 66
rect 6048 59 6090 61
rect 6146 59 6188 61
rect 6048 7 6060 59
rect 6176 7 6188 59
rect 6048 5 6090 7
rect 6146 5 6188 7
rect 6048 0 6188 5
rect 6216 0 6244 2272
rect 6272 66 6300 2338
rect 6328 2333 6468 2338
rect 6328 2331 6370 2333
rect 6426 2331 6468 2333
rect 6328 2279 6340 2331
rect 6456 2279 6468 2331
rect 6328 2277 6370 2279
rect 6426 2277 6468 2279
rect 6328 2272 6468 2277
rect 6328 94 6356 2272
rect 6384 66 6412 2244
rect 6272 61 6412 66
rect 6272 59 6314 61
rect 6370 59 6412 61
rect 6272 7 6284 59
rect 6400 7 6412 59
rect 6272 5 6314 7
rect 6370 5 6412 7
rect 6272 0 6412 5
rect 6440 0 6468 2272
rect 6496 66 6524 2338
rect 6552 2333 6692 2338
rect 6552 2331 6594 2333
rect 6650 2331 6692 2333
rect 6552 2279 6564 2331
rect 6680 2279 6692 2331
rect 6552 2277 6594 2279
rect 6650 2277 6692 2279
rect 6552 2272 6692 2277
rect 6552 94 6580 2272
rect 6608 66 6636 2244
rect 6496 61 6636 66
rect 6496 59 6538 61
rect 6594 59 6636 61
rect 6496 7 6508 59
rect 6624 7 6636 59
rect 6496 5 6538 7
rect 6594 5 6636 7
rect 6496 0 6636 5
rect 6664 0 6692 2272
rect 6720 66 6748 2338
rect 6776 2333 6916 2338
rect 6776 2331 6818 2333
rect 6874 2331 6916 2333
rect 6776 2279 6788 2331
rect 6904 2279 6916 2331
rect 6776 2277 6818 2279
rect 6874 2277 6916 2279
rect 6776 2272 6916 2277
rect 6776 94 6804 2272
rect 6832 66 6860 2244
rect 6720 61 6860 66
rect 6720 59 6762 61
rect 6818 59 6860 61
rect 6720 7 6732 59
rect 6848 7 6860 59
rect 6720 5 6762 7
rect 6818 5 6860 7
rect 6720 0 6860 5
rect 6888 0 6916 2272
rect 6944 66 6972 2338
rect 7000 2333 7140 2338
rect 7000 2331 7042 2333
rect 7098 2331 7140 2333
rect 7000 2279 7012 2331
rect 7128 2279 7140 2331
rect 7000 2277 7042 2279
rect 7098 2277 7140 2279
rect 7000 2272 7140 2277
rect 7000 94 7028 2272
rect 7056 66 7084 2244
rect 6944 61 7084 66
rect 6944 59 6986 61
rect 7042 59 7084 61
rect 6944 7 6956 59
rect 7072 7 7084 59
rect 6944 5 6986 7
rect 7042 5 7084 7
rect 6944 0 7084 5
rect 7112 0 7140 2272
rect 7168 66 7196 2338
rect 7224 2333 7364 2338
rect 7224 2331 7266 2333
rect 7322 2331 7364 2333
rect 7224 2279 7236 2331
rect 7352 2279 7364 2331
rect 7224 2277 7266 2279
rect 7322 2277 7364 2279
rect 7224 2272 7364 2277
rect 7224 94 7252 2272
rect 7280 66 7308 2244
rect 7168 61 7308 66
rect 7168 59 7210 61
rect 7266 59 7308 61
rect 7168 7 7180 59
rect 7296 7 7308 59
rect 7168 5 7210 7
rect 7266 5 7308 7
rect 7168 0 7308 5
rect 7336 0 7364 2272
rect 7392 66 7420 2338
rect 7448 2333 7588 2338
rect 7448 2331 7490 2333
rect 7546 2331 7588 2333
rect 7448 2279 7460 2331
rect 7576 2279 7588 2331
rect 7448 2277 7490 2279
rect 7546 2277 7588 2279
rect 7448 2272 7588 2277
rect 7448 94 7476 2272
rect 7504 66 7532 2244
rect 7392 61 7532 66
rect 7392 59 7434 61
rect 7490 59 7532 61
rect 7392 7 7404 59
rect 7520 7 7532 59
rect 7392 5 7434 7
rect 7490 5 7532 7
rect 7392 0 7532 5
rect 7560 0 7588 2272
rect 7616 66 7644 2338
rect 7672 2333 7812 2338
rect 7672 2331 7714 2333
rect 7770 2331 7812 2333
rect 7672 2279 7684 2331
rect 7800 2279 7812 2331
rect 7672 2277 7714 2279
rect 7770 2277 7812 2279
rect 7672 2272 7812 2277
rect 7672 94 7700 2272
rect 7728 66 7756 2244
rect 7616 61 7756 66
rect 7616 59 7658 61
rect 7714 59 7756 61
rect 7616 7 7628 59
rect 7744 7 7756 59
rect 7616 5 7658 7
rect 7714 5 7756 7
rect 7616 0 7756 5
rect 7784 0 7812 2272
rect 7840 66 7868 2338
rect 7896 2333 8036 2338
rect 7896 2331 7938 2333
rect 7994 2331 8036 2333
rect 7896 2279 7908 2331
rect 8024 2279 8036 2331
rect 7896 2277 7938 2279
rect 7994 2277 8036 2279
rect 7896 2272 8036 2277
rect 7896 94 7924 2272
rect 7952 66 7980 2244
rect 7840 61 7980 66
rect 7840 59 7882 61
rect 7938 59 7980 61
rect 7840 7 7852 59
rect 7968 7 7980 59
rect 7840 5 7882 7
rect 7938 5 7980 7
rect 7840 0 7980 5
rect 8008 0 8036 2272
rect 8064 66 8092 2338
rect 8120 2333 8260 2338
rect 8120 2331 8162 2333
rect 8218 2331 8260 2333
rect 8120 2279 8132 2331
rect 8248 2279 8260 2331
rect 8120 2277 8162 2279
rect 8218 2277 8260 2279
rect 8120 2272 8260 2277
rect 8120 94 8148 2272
rect 8176 66 8204 2244
rect 8064 61 8204 66
rect 8064 59 8106 61
rect 8162 59 8204 61
rect 8064 7 8076 59
rect 8192 7 8204 59
rect 8064 5 8106 7
rect 8162 5 8204 7
rect 8064 0 8204 5
rect 8232 0 8260 2272
rect 8288 66 8316 2338
rect 8344 2333 8484 2338
rect 8344 2331 8386 2333
rect 8442 2331 8484 2333
rect 8344 2279 8356 2331
rect 8472 2279 8484 2331
rect 8344 2277 8386 2279
rect 8442 2277 8484 2279
rect 8344 2272 8484 2277
rect 8344 94 8372 2272
rect 8400 66 8428 2244
rect 8288 61 8428 66
rect 8288 59 8330 61
rect 8386 59 8428 61
rect 8288 7 8300 59
rect 8416 7 8428 59
rect 8288 5 8330 7
rect 8386 5 8428 7
rect 8288 0 8428 5
rect 8456 0 8484 2272
rect 8512 66 8540 2338
rect 8568 2333 8708 2338
rect 8568 2331 8610 2333
rect 8666 2331 8708 2333
rect 8568 2279 8580 2331
rect 8696 2279 8708 2331
rect 8568 2277 8610 2279
rect 8666 2277 8708 2279
rect 8568 2272 8708 2277
rect 8568 94 8596 2272
rect 8624 66 8652 2244
rect 8512 61 8652 66
rect 8512 59 8554 61
rect 8610 59 8652 61
rect 8512 7 8524 59
rect 8640 7 8652 59
rect 8512 5 8554 7
rect 8610 5 8652 7
rect 8512 0 8652 5
rect 8680 0 8708 2272
rect 8736 66 8764 2338
rect 8792 2333 8932 2338
rect 8792 2331 8834 2333
rect 8890 2331 8932 2333
rect 8792 2279 8804 2331
rect 8920 2279 8932 2331
rect 8792 2277 8834 2279
rect 8890 2277 8932 2279
rect 8792 2272 8932 2277
rect 8792 94 8820 2272
rect 8848 66 8876 2244
rect 8736 61 8876 66
rect 8736 59 8778 61
rect 8834 59 8876 61
rect 8736 7 8748 59
rect 8864 7 8876 59
rect 8736 5 8778 7
rect 8834 5 8876 7
rect 8736 0 8876 5
rect 8904 0 8932 2272
rect 8960 66 8988 2338
rect 9016 2333 9156 2338
rect 9016 2331 9058 2333
rect 9114 2331 9156 2333
rect 9016 2279 9028 2331
rect 9144 2279 9156 2331
rect 9016 2277 9058 2279
rect 9114 2277 9156 2279
rect 9016 2272 9156 2277
rect 9016 94 9044 2272
rect 9072 66 9100 2244
rect 8960 61 9100 66
rect 8960 59 9002 61
rect 9058 59 9100 61
rect 8960 7 8972 59
rect 9088 7 9100 59
rect 8960 5 9002 7
rect 9058 5 9100 7
rect 8960 0 9100 5
rect 9128 0 9156 2272
rect 9184 66 9212 2338
rect 9240 2333 9380 2338
rect 9240 2331 9282 2333
rect 9338 2331 9380 2333
rect 9240 2279 9252 2331
rect 9368 2279 9380 2331
rect 9240 2277 9282 2279
rect 9338 2277 9380 2279
rect 9240 2272 9380 2277
rect 9240 94 9268 2272
rect 9296 66 9324 2244
rect 9184 61 9324 66
rect 9184 59 9226 61
rect 9282 59 9324 61
rect 9184 7 9196 59
rect 9312 7 9324 59
rect 9184 5 9226 7
rect 9282 5 9324 7
rect 9184 0 9324 5
rect 9352 0 9380 2272
rect 9408 66 9436 2338
rect 9464 2333 9604 2338
rect 9464 2331 9506 2333
rect 9562 2331 9604 2333
rect 9464 2279 9476 2331
rect 9592 2279 9604 2331
rect 9464 2277 9506 2279
rect 9562 2277 9604 2279
rect 9464 2272 9604 2277
rect 9464 94 9492 2272
rect 9520 66 9548 2244
rect 9408 61 9548 66
rect 9408 59 9450 61
rect 9506 59 9548 61
rect 9408 7 9420 59
rect 9536 7 9548 59
rect 9408 5 9450 7
rect 9506 5 9548 7
rect 9408 0 9548 5
rect 9576 0 9604 2272
rect 9632 66 9660 2338
rect 9688 2333 9828 2338
rect 9688 2331 9730 2333
rect 9786 2331 9828 2333
rect 9688 2279 9700 2331
rect 9816 2279 9828 2331
rect 9688 2277 9730 2279
rect 9786 2277 9828 2279
rect 9688 2272 9828 2277
rect 9688 94 9716 2272
rect 9744 66 9772 2244
rect 9632 61 9772 66
rect 9632 59 9674 61
rect 9730 59 9772 61
rect 9632 7 9644 59
rect 9760 7 9772 59
rect 9632 5 9674 7
rect 9730 5 9772 7
rect 9632 0 9772 5
rect 9800 0 9828 2272
rect 9856 66 9884 2338
rect 9912 2333 10052 2338
rect 9912 2331 9954 2333
rect 10010 2331 10052 2333
rect 9912 2279 9924 2331
rect 10040 2279 10052 2331
rect 9912 2277 9954 2279
rect 10010 2277 10052 2279
rect 9912 2272 10052 2277
rect 9912 94 9940 2272
rect 9968 66 9996 2244
rect 9856 61 9996 66
rect 9856 59 9898 61
rect 9954 59 9996 61
rect 9856 7 9868 59
rect 9984 7 9996 59
rect 9856 5 9898 7
rect 9954 5 9996 7
rect 9856 0 9996 5
rect 10024 0 10052 2272
rect 10080 66 10108 2338
rect 10136 2333 10276 2338
rect 10136 2331 10178 2333
rect 10234 2331 10276 2333
rect 10136 2279 10148 2331
rect 10264 2279 10276 2331
rect 10136 2277 10178 2279
rect 10234 2277 10276 2279
rect 10136 2272 10276 2277
rect 10136 94 10164 2272
rect 10192 66 10220 2244
rect 10080 61 10220 66
rect 10080 59 10122 61
rect 10178 59 10220 61
rect 10080 7 10092 59
rect 10208 7 10220 59
rect 10080 5 10122 7
rect 10178 5 10220 7
rect 10080 0 10220 5
rect 10248 0 10276 2272
rect 10304 66 10332 2338
rect 10360 2333 10500 2338
rect 10360 2331 10402 2333
rect 10458 2331 10500 2333
rect 10360 2279 10372 2331
rect 10488 2279 10500 2331
rect 10360 2277 10402 2279
rect 10458 2277 10500 2279
rect 10360 2272 10500 2277
rect 10360 94 10388 2272
rect 10416 66 10444 2244
rect 10304 61 10444 66
rect 10304 59 10346 61
rect 10402 59 10444 61
rect 10304 7 10316 59
rect 10432 7 10444 59
rect 10304 5 10346 7
rect 10402 5 10444 7
rect 10304 0 10444 5
rect 10472 0 10500 2272
rect 10528 66 10556 2338
rect 10584 2333 10724 2338
rect 10584 2331 10626 2333
rect 10682 2331 10724 2333
rect 10584 2279 10596 2331
rect 10712 2279 10724 2331
rect 10584 2277 10626 2279
rect 10682 2277 10724 2279
rect 10584 2272 10724 2277
rect 10584 94 10612 2272
rect 10640 66 10668 2244
rect 10528 61 10668 66
rect 10528 59 10570 61
rect 10626 59 10668 61
rect 10528 7 10540 59
rect 10656 7 10668 59
rect 10528 5 10570 7
rect 10626 5 10668 7
rect 10528 0 10668 5
rect 10696 0 10724 2272
rect 10752 66 10780 2338
rect 10808 2333 11146 2338
rect 10808 2331 10850 2333
rect 10906 2331 11146 2333
rect 10808 2279 10820 2331
rect 10936 2279 11146 2331
rect 10808 2277 10850 2279
rect 10906 2277 11146 2279
rect 10808 2272 11146 2277
rect 10808 94 10836 2272
rect 10864 66 10892 2244
rect 10752 61 10892 66
rect 10752 59 10794 61
rect 10850 59 10892 61
rect 10752 7 10764 59
rect 10880 7 10892 59
rect 10752 5 10794 7
rect 10850 5 10892 7
rect 10752 0 10892 5
rect 10920 0 10948 2272
rect 10976 66 11004 2244
rect 11032 94 11060 2272
rect 11088 66 11146 2244
rect 10976 61 11146 66
rect 10976 59 11018 61
rect 11074 59 11146 61
rect 10976 7 10988 59
rect 11104 7 11146 59
rect 10976 5 11018 7
rect 11074 5 11146 7
rect 10976 0 11146 5
<< via2 >>
rect 98 2331 154 2333
rect 98 2279 120 2331
rect 120 2279 132 2331
rect 132 2279 154 2331
rect 98 2277 154 2279
rect 42 59 98 61
rect 42 7 76 59
rect 76 7 88 59
rect 88 7 98 59
rect 42 5 98 7
rect 322 2331 378 2333
rect 322 2279 344 2331
rect 344 2279 356 2331
rect 356 2279 378 2331
rect 322 2277 378 2279
rect 266 59 322 61
rect 266 7 288 59
rect 288 7 300 59
rect 300 7 322 59
rect 266 5 322 7
rect 546 2331 602 2333
rect 546 2279 568 2331
rect 568 2279 580 2331
rect 580 2279 602 2331
rect 546 2277 602 2279
rect 490 59 546 61
rect 490 7 512 59
rect 512 7 524 59
rect 524 7 546 59
rect 490 5 546 7
rect 770 2331 826 2333
rect 770 2279 792 2331
rect 792 2279 804 2331
rect 804 2279 826 2331
rect 770 2277 826 2279
rect 714 59 770 61
rect 714 7 736 59
rect 736 7 748 59
rect 748 7 770 59
rect 714 5 770 7
rect 994 2331 1050 2333
rect 994 2279 1016 2331
rect 1016 2279 1028 2331
rect 1028 2279 1050 2331
rect 994 2277 1050 2279
rect 938 59 994 61
rect 938 7 960 59
rect 960 7 972 59
rect 972 7 994 59
rect 938 5 994 7
rect 1218 2331 1274 2333
rect 1218 2279 1240 2331
rect 1240 2279 1252 2331
rect 1252 2279 1274 2331
rect 1218 2277 1274 2279
rect 1162 59 1218 61
rect 1162 7 1184 59
rect 1184 7 1196 59
rect 1196 7 1218 59
rect 1162 5 1218 7
rect 1442 2331 1498 2333
rect 1442 2279 1464 2331
rect 1464 2279 1476 2331
rect 1476 2279 1498 2331
rect 1442 2277 1498 2279
rect 1386 59 1442 61
rect 1386 7 1408 59
rect 1408 7 1420 59
rect 1420 7 1442 59
rect 1386 5 1442 7
rect 1666 2331 1722 2333
rect 1666 2279 1688 2331
rect 1688 2279 1700 2331
rect 1700 2279 1722 2331
rect 1666 2277 1722 2279
rect 1610 59 1666 61
rect 1610 7 1632 59
rect 1632 7 1644 59
rect 1644 7 1666 59
rect 1610 5 1666 7
rect 1890 2331 1946 2333
rect 1890 2279 1912 2331
rect 1912 2279 1924 2331
rect 1924 2279 1946 2331
rect 1890 2277 1946 2279
rect 1834 59 1890 61
rect 1834 7 1856 59
rect 1856 7 1868 59
rect 1868 7 1890 59
rect 1834 5 1890 7
rect 2114 2331 2170 2333
rect 2114 2279 2136 2331
rect 2136 2279 2148 2331
rect 2148 2279 2170 2331
rect 2114 2277 2170 2279
rect 2058 59 2114 61
rect 2058 7 2080 59
rect 2080 7 2092 59
rect 2092 7 2114 59
rect 2058 5 2114 7
rect 2338 2331 2394 2333
rect 2338 2279 2360 2331
rect 2360 2279 2372 2331
rect 2372 2279 2394 2331
rect 2338 2277 2394 2279
rect 2282 59 2338 61
rect 2282 7 2304 59
rect 2304 7 2316 59
rect 2316 7 2338 59
rect 2282 5 2338 7
rect 2562 2331 2618 2333
rect 2562 2279 2584 2331
rect 2584 2279 2596 2331
rect 2596 2279 2618 2331
rect 2562 2277 2618 2279
rect 2506 59 2562 61
rect 2506 7 2528 59
rect 2528 7 2540 59
rect 2540 7 2562 59
rect 2506 5 2562 7
rect 2786 2331 2842 2333
rect 2786 2279 2808 2331
rect 2808 2279 2820 2331
rect 2820 2279 2842 2331
rect 2786 2277 2842 2279
rect 2730 59 2786 61
rect 2730 7 2752 59
rect 2752 7 2764 59
rect 2764 7 2786 59
rect 2730 5 2786 7
rect 3010 2331 3066 2333
rect 3010 2279 3032 2331
rect 3032 2279 3044 2331
rect 3044 2279 3066 2331
rect 3010 2277 3066 2279
rect 2954 59 3010 61
rect 2954 7 2976 59
rect 2976 7 2988 59
rect 2988 7 3010 59
rect 2954 5 3010 7
rect 3234 2331 3290 2333
rect 3234 2279 3256 2331
rect 3256 2279 3268 2331
rect 3268 2279 3290 2331
rect 3234 2277 3290 2279
rect 3178 59 3234 61
rect 3178 7 3200 59
rect 3200 7 3212 59
rect 3212 7 3234 59
rect 3178 5 3234 7
rect 3458 2331 3514 2333
rect 3458 2279 3480 2331
rect 3480 2279 3492 2331
rect 3492 2279 3514 2331
rect 3458 2277 3514 2279
rect 3402 59 3458 61
rect 3402 7 3424 59
rect 3424 7 3436 59
rect 3436 7 3458 59
rect 3402 5 3458 7
rect 3682 2331 3738 2333
rect 3682 2279 3704 2331
rect 3704 2279 3716 2331
rect 3716 2279 3738 2331
rect 3682 2277 3738 2279
rect 3626 59 3682 61
rect 3626 7 3648 59
rect 3648 7 3660 59
rect 3660 7 3682 59
rect 3626 5 3682 7
rect 3906 2331 3962 2333
rect 3906 2279 3928 2331
rect 3928 2279 3940 2331
rect 3940 2279 3962 2331
rect 3906 2277 3962 2279
rect 3850 59 3906 61
rect 3850 7 3872 59
rect 3872 7 3884 59
rect 3884 7 3906 59
rect 3850 5 3906 7
rect 4130 2331 4186 2333
rect 4130 2279 4152 2331
rect 4152 2279 4164 2331
rect 4164 2279 4186 2331
rect 4130 2277 4186 2279
rect 4074 59 4130 61
rect 4074 7 4096 59
rect 4096 7 4108 59
rect 4108 7 4130 59
rect 4074 5 4130 7
rect 4354 2331 4410 2333
rect 4354 2279 4376 2331
rect 4376 2279 4388 2331
rect 4388 2279 4410 2331
rect 4354 2277 4410 2279
rect 4298 59 4354 61
rect 4298 7 4320 59
rect 4320 7 4332 59
rect 4332 7 4354 59
rect 4298 5 4354 7
rect 4578 2331 4634 2333
rect 4578 2279 4600 2331
rect 4600 2279 4612 2331
rect 4612 2279 4634 2331
rect 4578 2277 4634 2279
rect 4522 59 4578 61
rect 4522 7 4544 59
rect 4544 7 4556 59
rect 4556 7 4578 59
rect 4522 5 4578 7
rect 4802 2331 4858 2333
rect 4802 2279 4824 2331
rect 4824 2279 4836 2331
rect 4836 2279 4858 2331
rect 4802 2277 4858 2279
rect 4746 59 4802 61
rect 4746 7 4768 59
rect 4768 7 4780 59
rect 4780 7 4802 59
rect 4746 5 4802 7
rect 5026 2331 5082 2333
rect 5026 2279 5048 2331
rect 5048 2279 5060 2331
rect 5060 2279 5082 2331
rect 5026 2277 5082 2279
rect 4970 59 5026 61
rect 4970 7 4992 59
rect 4992 7 5004 59
rect 5004 7 5026 59
rect 4970 5 5026 7
rect 5250 2331 5306 2333
rect 5250 2279 5272 2331
rect 5272 2279 5284 2331
rect 5284 2279 5306 2331
rect 5250 2277 5306 2279
rect 5194 59 5250 61
rect 5194 7 5216 59
rect 5216 7 5228 59
rect 5228 7 5250 59
rect 5194 5 5250 7
rect 5474 2331 5530 2333
rect 5474 2279 5496 2331
rect 5496 2279 5508 2331
rect 5508 2279 5530 2331
rect 5474 2277 5530 2279
rect 5418 59 5474 61
rect 5418 7 5440 59
rect 5440 7 5452 59
rect 5452 7 5474 59
rect 5418 5 5474 7
rect 5698 2331 5754 2333
rect 5698 2279 5720 2331
rect 5720 2279 5732 2331
rect 5732 2279 5754 2331
rect 5698 2277 5754 2279
rect 5642 59 5698 61
rect 5642 7 5664 59
rect 5664 7 5676 59
rect 5676 7 5698 59
rect 5642 5 5698 7
rect 5922 2331 5978 2333
rect 5922 2279 5944 2331
rect 5944 2279 5956 2331
rect 5956 2279 5978 2331
rect 5922 2277 5978 2279
rect 5866 59 5922 61
rect 5866 7 5888 59
rect 5888 7 5900 59
rect 5900 7 5922 59
rect 5866 5 5922 7
rect 6146 2331 6202 2333
rect 6146 2279 6168 2331
rect 6168 2279 6180 2331
rect 6180 2279 6202 2331
rect 6146 2277 6202 2279
rect 6090 59 6146 61
rect 6090 7 6112 59
rect 6112 7 6124 59
rect 6124 7 6146 59
rect 6090 5 6146 7
rect 6370 2331 6426 2333
rect 6370 2279 6392 2331
rect 6392 2279 6404 2331
rect 6404 2279 6426 2331
rect 6370 2277 6426 2279
rect 6314 59 6370 61
rect 6314 7 6336 59
rect 6336 7 6348 59
rect 6348 7 6370 59
rect 6314 5 6370 7
rect 6594 2331 6650 2333
rect 6594 2279 6616 2331
rect 6616 2279 6628 2331
rect 6628 2279 6650 2331
rect 6594 2277 6650 2279
rect 6538 59 6594 61
rect 6538 7 6560 59
rect 6560 7 6572 59
rect 6572 7 6594 59
rect 6538 5 6594 7
rect 6818 2331 6874 2333
rect 6818 2279 6840 2331
rect 6840 2279 6852 2331
rect 6852 2279 6874 2331
rect 6818 2277 6874 2279
rect 6762 59 6818 61
rect 6762 7 6784 59
rect 6784 7 6796 59
rect 6796 7 6818 59
rect 6762 5 6818 7
rect 7042 2331 7098 2333
rect 7042 2279 7064 2331
rect 7064 2279 7076 2331
rect 7076 2279 7098 2331
rect 7042 2277 7098 2279
rect 6986 59 7042 61
rect 6986 7 7008 59
rect 7008 7 7020 59
rect 7020 7 7042 59
rect 6986 5 7042 7
rect 7266 2331 7322 2333
rect 7266 2279 7288 2331
rect 7288 2279 7300 2331
rect 7300 2279 7322 2331
rect 7266 2277 7322 2279
rect 7210 59 7266 61
rect 7210 7 7232 59
rect 7232 7 7244 59
rect 7244 7 7266 59
rect 7210 5 7266 7
rect 7490 2331 7546 2333
rect 7490 2279 7512 2331
rect 7512 2279 7524 2331
rect 7524 2279 7546 2331
rect 7490 2277 7546 2279
rect 7434 59 7490 61
rect 7434 7 7456 59
rect 7456 7 7468 59
rect 7468 7 7490 59
rect 7434 5 7490 7
rect 7714 2331 7770 2333
rect 7714 2279 7736 2331
rect 7736 2279 7748 2331
rect 7748 2279 7770 2331
rect 7714 2277 7770 2279
rect 7658 59 7714 61
rect 7658 7 7680 59
rect 7680 7 7692 59
rect 7692 7 7714 59
rect 7658 5 7714 7
rect 7938 2331 7994 2333
rect 7938 2279 7960 2331
rect 7960 2279 7972 2331
rect 7972 2279 7994 2331
rect 7938 2277 7994 2279
rect 7882 59 7938 61
rect 7882 7 7904 59
rect 7904 7 7916 59
rect 7916 7 7938 59
rect 7882 5 7938 7
rect 8162 2331 8218 2333
rect 8162 2279 8184 2331
rect 8184 2279 8196 2331
rect 8196 2279 8218 2331
rect 8162 2277 8218 2279
rect 8106 59 8162 61
rect 8106 7 8128 59
rect 8128 7 8140 59
rect 8140 7 8162 59
rect 8106 5 8162 7
rect 8386 2331 8442 2333
rect 8386 2279 8408 2331
rect 8408 2279 8420 2331
rect 8420 2279 8442 2331
rect 8386 2277 8442 2279
rect 8330 59 8386 61
rect 8330 7 8352 59
rect 8352 7 8364 59
rect 8364 7 8386 59
rect 8330 5 8386 7
rect 8610 2331 8666 2333
rect 8610 2279 8632 2331
rect 8632 2279 8644 2331
rect 8644 2279 8666 2331
rect 8610 2277 8666 2279
rect 8554 59 8610 61
rect 8554 7 8576 59
rect 8576 7 8588 59
rect 8588 7 8610 59
rect 8554 5 8610 7
rect 8834 2331 8890 2333
rect 8834 2279 8856 2331
rect 8856 2279 8868 2331
rect 8868 2279 8890 2331
rect 8834 2277 8890 2279
rect 8778 59 8834 61
rect 8778 7 8800 59
rect 8800 7 8812 59
rect 8812 7 8834 59
rect 8778 5 8834 7
rect 9058 2331 9114 2333
rect 9058 2279 9080 2331
rect 9080 2279 9092 2331
rect 9092 2279 9114 2331
rect 9058 2277 9114 2279
rect 9002 59 9058 61
rect 9002 7 9024 59
rect 9024 7 9036 59
rect 9036 7 9058 59
rect 9002 5 9058 7
rect 9282 2331 9338 2333
rect 9282 2279 9304 2331
rect 9304 2279 9316 2331
rect 9316 2279 9338 2331
rect 9282 2277 9338 2279
rect 9226 59 9282 61
rect 9226 7 9248 59
rect 9248 7 9260 59
rect 9260 7 9282 59
rect 9226 5 9282 7
rect 9506 2331 9562 2333
rect 9506 2279 9528 2331
rect 9528 2279 9540 2331
rect 9540 2279 9562 2331
rect 9506 2277 9562 2279
rect 9450 59 9506 61
rect 9450 7 9472 59
rect 9472 7 9484 59
rect 9484 7 9506 59
rect 9450 5 9506 7
rect 9730 2331 9786 2333
rect 9730 2279 9752 2331
rect 9752 2279 9764 2331
rect 9764 2279 9786 2331
rect 9730 2277 9786 2279
rect 9674 59 9730 61
rect 9674 7 9696 59
rect 9696 7 9708 59
rect 9708 7 9730 59
rect 9674 5 9730 7
rect 9954 2331 10010 2333
rect 9954 2279 9976 2331
rect 9976 2279 9988 2331
rect 9988 2279 10010 2331
rect 9954 2277 10010 2279
rect 9898 59 9954 61
rect 9898 7 9920 59
rect 9920 7 9932 59
rect 9932 7 9954 59
rect 9898 5 9954 7
rect 10178 2331 10234 2333
rect 10178 2279 10200 2331
rect 10200 2279 10212 2331
rect 10212 2279 10234 2331
rect 10178 2277 10234 2279
rect 10122 59 10178 61
rect 10122 7 10144 59
rect 10144 7 10156 59
rect 10156 7 10178 59
rect 10122 5 10178 7
rect 10402 2331 10458 2333
rect 10402 2279 10424 2331
rect 10424 2279 10436 2331
rect 10436 2279 10458 2331
rect 10402 2277 10458 2279
rect 10346 59 10402 61
rect 10346 7 10368 59
rect 10368 7 10380 59
rect 10380 7 10402 59
rect 10346 5 10402 7
rect 10626 2331 10682 2333
rect 10626 2279 10648 2331
rect 10648 2279 10660 2331
rect 10660 2279 10682 2331
rect 10626 2277 10682 2279
rect 10570 59 10626 61
rect 10570 7 10592 59
rect 10592 7 10604 59
rect 10604 7 10626 59
rect 10570 5 10626 7
rect 10850 2331 10906 2333
rect 10850 2279 10872 2331
rect 10872 2279 10884 2331
rect 10884 2279 10906 2331
rect 10850 2277 10906 2279
rect 10794 59 10850 61
rect 10794 7 10816 59
rect 10816 7 10828 59
rect 10828 7 10850 59
rect 10794 5 10850 7
rect 11018 59 11074 61
rect 11018 7 11040 59
rect 11040 7 11052 59
rect 11052 7 11074 59
rect 11018 5 11074 7
<< metal3 >>
rect 0 2337 11146 2338
rect 0 2273 28 2337
rect 92 2333 108 2337
rect 92 2277 98 2333
rect 92 2273 108 2277
rect 172 2273 188 2337
rect 252 2273 268 2337
rect 332 2333 348 2337
rect 332 2273 348 2277
rect 412 2273 428 2337
rect 492 2273 508 2337
rect 572 2333 588 2337
rect 572 2273 588 2277
rect 652 2273 668 2337
rect 732 2273 748 2337
rect 812 2333 828 2337
rect 826 2277 828 2333
rect 812 2273 828 2277
rect 892 2273 908 2337
rect 972 2273 988 2337
rect 1052 2273 1068 2337
rect 1132 2273 1148 2337
rect 1212 2333 1228 2337
rect 1212 2277 1218 2333
rect 1212 2273 1228 2277
rect 1292 2273 1308 2337
rect 1372 2273 1388 2337
rect 1452 2333 1468 2337
rect 1452 2273 1468 2277
rect 1532 2273 1548 2337
rect 1612 2273 1628 2337
rect 1692 2333 1708 2337
rect 1692 2273 1708 2277
rect 1772 2273 1788 2337
rect 1852 2273 1868 2337
rect 1932 2333 1948 2337
rect 1946 2277 1948 2333
rect 1932 2273 1948 2277
rect 2012 2273 2028 2337
rect 2092 2273 2108 2337
rect 2172 2273 2188 2337
rect 2252 2273 2268 2337
rect 2332 2333 2348 2337
rect 2332 2277 2338 2333
rect 2332 2273 2348 2277
rect 2412 2273 2428 2337
rect 2492 2273 2508 2337
rect 2572 2333 2588 2337
rect 2572 2273 2588 2277
rect 2652 2273 2668 2337
rect 2732 2273 2748 2337
rect 2812 2333 2828 2337
rect 2812 2273 2828 2277
rect 2892 2273 2908 2337
rect 2972 2273 2988 2337
rect 3052 2333 3068 2337
rect 3066 2277 3068 2333
rect 3052 2273 3068 2277
rect 3132 2273 3148 2337
rect 3212 2273 3228 2337
rect 3292 2273 3308 2337
rect 3372 2273 3388 2337
rect 3452 2333 3468 2337
rect 3452 2277 3458 2333
rect 3452 2273 3468 2277
rect 3532 2273 3548 2337
rect 3612 2273 3628 2337
rect 3692 2333 3708 2337
rect 3692 2273 3708 2277
rect 3772 2273 3788 2337
rect 3852 2273 3868 2337
rect 3932 2333 3948 2337
rect 3932 2273 3948 2277
rect 4012 2273 4028 2337
rect 4092 2273 4108 2337
rect 4172 2333 4188 2337
rect 4186 2277 4188 2333
rect 4172 2273 4188 2277
rect 4252 2273 4268 2337
rect 4332 2273 4348 2337
rect 4412 2273 4428 2337
rect 4492 2273 4508 2337
rect 4572 2333 4588 2337
rect 4572 2277 4578 2333
rect 4572 2273 4588 2277
rect 4652 2273 4668 2337
rect 4732 2273 4748 2337
rect 4812 2333 4828 2337
rect 4812 2273 4828 2277
rect 4892 2273 4908 2337
rect 4972 2273 4988 2337
rect 5052 2333 5068 2337
rect 5052 2273 5068 2277
rect 5132 2273 5148 2337
rect 5212 2273 5228 2337
rect 5292 2333 5308 2337
rect 5306 2277 5308 2333
rect 5292 2273 5308 2277
rect 5372 2273 5388 2337
rect 5452 2273 5468 2337
rect 5532 2273 5548 2337
rect 5612 2273 5628 2337
rect 5692 2333 5708 2337
rect 5692 2277 5698 2333
rect 5692 2273 5708 2277
rect 5772 2273 5788 2337
rect 5852 2273 5868 2337
rect 5932 2333 5948 2337
rect 5932 2273 5948 2277
rect 6012 2273 6028 2337
rect 6092 2273 6108 2337
rect 6172 2333 6188 2337
rect 6172 2273 6188 2277
rect 6252 2273 6268 2337
rect 6332 2273 6348 2337
rect 6412 2333 6428 2337
rect 6426 2277 6428 2333
rect 6412 2273 6428 2277
rect 6492 2273 6508 2337
rect 6572 2273 6588 2337
rect 6652 2273 6668 2337
rect 6732 2273 6748 2337
rect 6812 2333 6828 2337
rect 6812 2277 6818 2333
rect 6812 2273 6828 2277
rect 6892 2273 6908 2337
rect 6972 2273 6988 2337
rect 7052 2333 7068 2337
rect 7052 2273 7068 2277
rect 7132 2273 7148 2337
rect 7212 2273 7228 2337
rect 7292 2333 7308 2337
rect 7292 2273 7308 2277
rect 7372 2273 7388 2337
rect 7452 2273 7468 2337
rect 7532 2333 7548 2337
rect 7546 2277 7548 2333
rect 7532 2273 7548 2277
rect 7612 2273 7628 2337
rect 7692 2273 7708 2337
rect 7772 2273 7788 2337
rect 7852 2273 7868 2337
rect 7932 2333 7948 2337
rect 7932 2277 7938 2333
rect 7932 2273 7948 2277
rect 8012 2273 8028 2337
rect 8092 2273 8108 2337
rect 8172 2333 8188 2337
rect 8172 2273 8188 2277
rect 8252 2273 8268 2337
rect 8332 2273 8348 2337
rect 8412 2333 8428 2337
rect 8412 2273 8428 2277
rect 8492 2273 8508 2337
rect 8572 2273 8588 2337
rect 8652 2333 8668 2337
rect 8666 2277 8668 2333
rect 8652 2273 8668 2277
rect 8732 2273 8748 2337
rect 8812 2273 8828 2337
rect 8892 2273 8908 2337
rect 8972 2273 8988 2337
rect 9052 2333 9068 2337
rect 9052 2277 9058 2333
rect 9052 2273 9068 2277
rect 9132 2273 9148 2337
rect 9212 2273 9228 2337
rect 9292 2333 9308 2337
rect 9292 2273 9308 2277
rect 9372 2273 9388 2337
rect 9452 2273 9468 2337
rect 9532 2333 9548 2337
rect 9532 2273 9548 2277
rect 9612 2273 9628 2337
rect 9692 2273 9708 2337
rect 9772 2333 9788 2337
rect 9786 2277 9788 2333
rect 9772 2273 9788 2277
rect 9852 2273 9868 2337
rect 9932 2273 9948 2337
rect 10012 2273 10028 2337
rect 10092 2273 10108 2337
rect 10172 2333 10188 2337
rect 10172 2277 10178 2333
rect 10172 2273 10188 2277
rect 10252 2273 10268 2337
rect 10332 2273 10348 2337
rect 10412 2333 10428 2337
rect 10412 2273 10428 2277
rect 10492 2273 10508 2337
rect 10572 2273 10588 2337
rect 10652 2333 10668 2337
rect 10652 2273 10668 2277
rect 10732 2273 10748 2337
rect 10812 2273 10828 2337
rect 10892 2333 10908 2337
rect 10906 2277 10908 2333
rect 10892 2273 10908 2277
rect 10972 2273 10988 2337
rect 11052 2273 11146 2337
rect 0 2272 11146 2273
rect 0 126 60 2272
rect 120 66 180 2212
rect 240 126 300 2272
rect 360 66 420 2212
rect 480 126 540 2272
rect 600 66 660 2212
rect 720 126 780 2272
rect 840 66 900 2212
rect 960 126 1020 2272
rect 1080 66 1140 2212
rect 1200 126 1260 2272
rect 1320 66 1380 2212
rect 1440 126 1500 2272
rect 1560 66 1620 2212
rect 1680 126 1740 2272
rect 1800 66 1860 2212
rect 1920 126 1980 2272
rect 2040 66 2100 2212
rect 2160 126 2220 2272
rect 2280 66 2340 2212
rect 2400 126 2460 2272
rect 2520 66 2580 2212
rect 2640 126 2700 2272
rect 2760 66 2820 2212
rect 2880 126 2940 2272
rect 3000 66 3060 2212
rect 3120 126 3180 2272
rect 3240 66 3300 2212
rect 3360 126 3420 2272
rect 3480 66 3540 2212
rect 3600 126 3660 2272
rect 3720 66 3780 2212
rect 3840 126 3900 2272
rect 3960 66 4020 2212
rect 4080 126 4140 2272
rect 4200 66 4260 2212
rect 4320 126 4380 2272
rect 4440 66 4500 2212
rect 4560 126 4620 2272
rect 4680 66 4740 2212
rect 4800 126 4860 2272
rect 4920 66 4980 2212
rect 5040 126 5100 2272
rect 5160 66 5220 2212
rect 5280 126 5340 2272
rect 5400 66 5460 2212
rect 5520 126 5580 2272
rect 5640 66 5700 2212
rect 5760 126 5820 2272
rect 5880 66 5940 2212
rect 6000 126 6060 2272
rect 6120 66 6180 2212
rect 6240 126 6300 2272
rect 6360 66 6420 2212
rect 6480 126 6540 2272
rect 6600 66 6660 2212
rect 6720 126 6780 2272
rect 6840 66 6900 2212
rect 6960 126 7020 2272
rect 7080 66 7140 2212
rect 7200 126 7260 2272
rect 7320 66 7380 2212
rect 7440 126 7500 2272
rect 7560 66 7620 2212
rect 7680 126 7740 2272
rect 7800 66 7860 2212
rect 7920 126 7980 2272
rect 8040 66 8100 2212
rect 8160 126 8220 2272
rect 8280 66 8340 2212
rect 8400 126 8460 2272
rect 8520 66 8580 2212
rect 8640 126 8700 2272
rect 8760 66 8820 2212
rect 8880 126 8940 2272
rect 9000 66 9060 2212
rect 9120 126 9180 2272
rect 9240 66 9300 2212
rect 9360 126 9420 2272
rect 9480 66 9540 2212
rect 9600 126 9660 2272
rect 9720 66 9780 2212
rect 9840 126 9900 2272
rect 9960 66 10020 2212
rect 10080 126 10140 2272
rect 10200 66 10260 2212
rect 10320 126 10380 2272
rect 10440 66 10500 2212
rect 10560 126 10620 2272
rect 10680 66 10740 2212
rect 10800 126 10860 2272
rect 10920 66 10980 2212
rect 11040 126 11146 2272
rect 0 65 11146 66
rect 0 1 28 65
rect 92 61 108 65
rect 98 5 108 61
rect 92 1 108 5
rect 172 1 188 65
rect 252 61 268 65
rect 252 5 266 61
rect 252 1 268 5
rect 332 1 348 65
rect 412 1 428 65
rect 492 61 508 65
rect 492 1 508 5
rect 572 1 588 65
rect 652 1 668 65
rect 732 61 748 65
rect 732 1 748 5
rect 812 1 828 65
rect 892 1 908 65
rect 972 61 988 65
rect 972 1 988 5
rect 1052 1 1068 65
rect 1132 1 1148 65
rect 1212 61 1228 65
rect 1218 5 1228 61
rect 1212 1 1228 5
rect 1292 1 1308 65
rect 1372 61 1388 65
rect 1372 5 1386 61
rect 1372 1 1388 5
rect 1452 1 1468 65
rect 1532 1 1548 65
rect 1612 61 1628 65
rect 1612 1 1628 5
rect 1692 1 1708 65
rect 1772 1 1788 65
rect 1852 61 1868 65
rect 1852 1 1868 5
rect 1932 1 1948 65
rect 2012 1 2028 65
rect 2092 61 2108 65
rect 2092 1 2108 5
rect 2172 1 2188 65
rect 2252 1 2268 65
rect 2332 61 2348 65
rect 2338 5 2348 61
rect 2332 1 2348 5
rect 2412 1 2428 65
rect 2492 61 2508 65
rect 2492 5 2506 61
rect 2492 1 2508 5
rect 2572 1 2588 65
rect 2652 1 2668 65
rect 2732 61 2748 65
rect 2732 1 2748 5
rect 2812 1 2828 65
rect 2892 1 2908 65
rect 2972 61 2988 65
rect 2972 1 2988 5
rect 3052 1 3068 65
rect 3132 1 3148 65
rect 3212 61 3228 65
rect 3212 1 3228 5
rect 3292 1 3308 65
rect 3372 1 3388 65
rect 3452 61 3468 65
rect 3458 5 3468 61
rect 3452 1 3468 5
rect 3532 1 3548 65
rect 3612 61 3628 65
rect 3612 5 3626 61
rect 3612 1 3628 5
rect 3692 1 3708 65
rect 3772 1 3788 65
rect 3852 61 3868 65
rect 3852 1 3868 5
rect 3932 1 3948 65
rect 4012 1 4028 65
rect 4092 61 4108 65
rect 4092 1 4108 5
rect 4172 1 4188 65
rect 4252 1 4268 65
rect 4332 61 4348 65
rect 4332 1 4348 5
rect 4412 1 4428 65
rect 4492 1 4508 65
rect 4572 61 4588 65
rect 4578 5 4588 61
rect 4572 1 4588 5
rect 4652 1 4668 65
rect 4732 61 4748 65
rect 4732 5 4746 61
rect 4732 1 4748 5
rect 4812 1 4828 65
rect 4892 1 4908 65
rect 4972 61 4988 65
rect 4972 1 4988 5
rect 5052 1 5068 65
rect 5132 1 5148 65
rect 5212 61 5228 65
rect 5212 1 5228 5
rect 5292 1 5308 65
rect 5372 1 5388 65
rect 5452 61 5468 65
rect 5452 1 5468 5
rect 5532 1 5548 65
rect 5612 1 5628 65
rect 5692 61 5708 65
rect 5698 5 5708 61
rect 5692 1 5708 5
rect 5772 1 5788 65
rect 5852 61 5868 65
rect 5852 5 5866 61
rect 5852 1 5868 5
rect 5932 1 5948 65
rect 6012 1 6028 65
rect 6092 61 6108 65
rect 6092 1 6108 5
rect 6172 1 6188 65
rect 6252 1 6268 65
rect 6332 61 6348 65
rect 6332 1 6348 5
rect 6412 1 6428 65
rect 6492 1 6508 65
rect 6572 61 6588 65
rect 6572 1 6588 5
rect 6652 1 6668 65
rect 6732 1 6748 65
rect 6812 61 6828 65
rect 6818 5 6828 61
rect 6812 1 6828 5
rect 6892 1 6908 65
rect 6972 61 6988 65
rect 6972 5 6986 61
rect 6972 1 6988 5
rect 7052 1 7068 65
rect 7132 1 7148 65
rect 7212 61 7228 65
rect 7212 1 7228 5
rect 7292 1 7308 65
rect 7372 1 7388 65
rect 7452 61 7468 65
rect 7452 1 7468 5
rect 7532 1 7548 65
rect 7612 1 7628 65
rect 7692 61 7708 65
rect 7692 1 7708 5
rect 7772 1 7788 65
rect 7852 1 7868 65
rect 7932 61 7948 65
rect 7938 5 7948 61
rect 7932 1 7948 5
rect 8012 1 8028 65
rect 8092 61 8108 65
rect 8092 5 8106 61
rect 8092 1 8108 5
rect 8172 1 8188 65
rect 8252 1 8268 65
rect 8332 61 8348 65
rect 8332 1 8348 5
rect 8412 1 8428 65
rect 8492 1 8508 65
rect 8572 61 8588 65
rect 8572 1 8588 5
rect 8652 1 8668 65
rect 8732 1 8748 65
rect 8812 61 8828 65
rect 8812 1 8828 5
rect 8892 1 8908 65
rect 8972 1 8988 65
rect 9052 61 9068 65
rect 9058 5 9068 61
rect 9052 1 9068 5
rect 9132 1 9148 65
rect 9212 61 9228 65
rect 9212 5 9226 61
rect 9212 1 9228 5
rect 9292 1 9308 65
rect 9372 1 9388 65
rect 9452 61 9468 65
rect 9452 1 9468 5
rect 9532 1 9548 65
rect 9612 1 9628 65
rect 9692 61 9708 65
rect 9692 1 9708 5
rect 9772 1 9788 65
rect 9852 1 9868 65
rect 9932 61 9948 65
rect 9932 1 9948 5
rect 10012 1 10028 65
rect 10092 1 10108 65
rect 10172 61 10188 65
rect 10178 5 10188 61
rect 10172 1 10188 5
rect 10252 1 10268 65
rect 10332 61 10348 65
rect 10332 5 10346 61
rect 10332 1 10348 5
rect 10412 1 10428 65
rect 10492 1 10508 65
rect 10572 61 10588 65
rect 10572 1 10588 5
rect 10652 1 10668 65
rect 10732 1 10748 65
rect 10812 61 10828 65
rect 10812 1 10828 5
rect 10892 1 10908 65
rect 10972 1 10988 65
rect 11052 61 11146 65
rect 11074 5 11146 61
rect 11052 1 11146 5
rect 0 0 11146 1
<< via3 >>
rect 28 2273 92 2337
rect 108 2333 172 2337
rect 108 2277 154 2333
rect 154 2277 172 2333
rect 108 2273 172 2277
rect 188 2273 252 2337
rect 268 2333 332 2337
rect 348 2333 412 2337
rect 268 2277 322 2333
rect 322 2277 332 2333
rect 348 2277 378 2333
rect 378 2277 412 2333
rect 268 2273 332 2277
rect 348 2273 412 2277
rect 428 2273 492 2337
rect 508 2333 572 2337
rect 588 2333 652 2337
rect 508 2277 546 2333
rect 546 2277 572 2333
rect 588 2277 602 2333
rect 602 2277 652 2333
rect 508 2273 572 2277
rect 588 2273 652 2277
rect 668 2273 732 2337
rect 748 2333 812 2337
rect 748 2277 770 2333
rect 770 2277 812 2333
rect 748 2273 812 2277
rect 828 2273 892 2337
rect 908 2273 972 2337
rect 988 2333 1052 2337
rect 988 2277 994 2333
rect 994 2277 1050 2333
rect 1050 2277 1052 2333
rect 988 2273 1052 2277
rect 1068 2273 1132 2337
rect 1148 2273 1212 2337
rect 1228 2333 1292 2337
rect 1228 2277 1274 2333
rect 1274 2277 1292 2333
rect 1228 2273 1292 2277
rect 1308 2273 1372 2337
rect 1388 2333 1452 2337
rect 1468 2333 1532 2337
rect 1388 2277 1442 2333
rect 1442 2277 1452 2333
rect 1468 2277 1498 2333
rect 1498 2277 1532 2333
rect 1388 2273 1452 2277
rect 1468 2273 1532 2277
rect 1548 2273 1612 2337
rect 1628 2333 1692 2337
rect 1708 2333 1772 2337
rect 1628 2277 1666 2333
rect 1666 2277 1692 2333
rect 1708 2277 1722 2333
rect 1722 2277 1772 2333
rect 1628 2273 1692 2277
rect 1708 2273 1772 2277
rect 1788 2273 1852 2337
rect 1868 2333 1932 2337
rect 1868 2277 1890 2333
rect 1890 2277 1932 2333
rect 1868 2273 1932 2277
rect 1948 2273 2012 2337
rect 2028 2273 2092 2337
rect 2108 2333 2172 2337
rect 2108 2277 2114 2333
rect 2114 2277 2170 2333
rect 2170 2277 2172 2333
rect 2108 2273 2172 2277
rect 2188 2273 2252 2337
rect 2268 2273 2332 2337
rect 2348 2333 2412 2337
rect 2348 2277 2394 2333
rect 2394 2277 2412 2333
rect 2348 2273 2412 2277
rect 2428 2273 2492 2337
rect 2508 2333 2572 2337
rect 2588 2333 2652 2337
rect 2508 2277 2562 2333
rect 2562 2277 2572 2333
rect 2588 2277 2618 2333
rect 2618 2277 2652 2333
rect 2508 2273 2572 2277
rect 2588 2273 2652 2277
rect 2668 2273 2732 2337
rect 2748 2333 2812 2337
rect 2828 2333 2892 2337
rect 2748 2277 2786 2333
rect 2786 2277 2812 2333
rect 2828 2277 2842 2333
rect 2842 2277 2892 2333
rect 2748 2273 2812 2277
rect 2828 2273 2892 2277
rect 2908 2273 2972 2337
rect 2988 2333 3052 2337
rect 2988 2277 3010 2333
rect 3010 2277 3052 2333
rect 2988 2273 3052 2277
rect 3068 2273 3132 2337
rect 3148 2273 3212 2337
rect 3228 2333 3292 2337
rect 3228 2277 3234 2333
rect 3234 2277 3290 2333
rect 3290 2277 3292 2333
rect 3228 2273 3292 2277
rect 3308 2273 3372 2337
rect 3388 2273 3452 2337
rect 3468 2333 3532 2337
rect 3468 2277 3514 2333
rect 3514 2277 3532 2333
rect 3468 2273 3532 2277
rect 3548 2273 3612 2337
rect 3628 2333 3692 2337
rect 3708 2333 3772 2337
rect 3628 2277 3682 2333
rect 3682 2277 3692 2333
rect 3708 2277 3738 2333
rect 3738 2277 3772 2333
rect 3628 2273 3692 2277
rect 3708 2273 3772 2277
rect 3788 2273 3852 2337
rect 3868 2333 3932 2337
rect 3948 2333 4012 2337
rect 3868 2277 3906 2333
rect 3906 2277 3932 2333
rect 3948 2277 3962 2333
rect 3962 2277 4012 2333
rect 3868 2273 3932 2277
rect 3948 2273 4012 2277
rect 4028 2273 4092 2337
rect 4108 2333 4172 2337
rect 4108 2277 4130 2333
rect 4130 2277 4172 2333
rect 4108 2273 4172 2277
rect 4188 2273 4252 2337
rect 4268 2273 4332 2337
rect 4348 2333 4412 2337
rect 4348 2277 4354 2333
rect 4354 2277 4410 2333
rect 4410 2277 4412 2333
rect 4348 2273 4412 2277
rect 4428 2273 4492 2337
rect 4508 2273 4572 2337
rect 4588 2333 4652 2337
rect 4588 2277 4634 2333
rect 4634 2277 4652 2333
rect 4588 2273 4652 2277
rect 4668 2273 4732 2337
rect 4748 2333 4812 2337
rect 4828 2333 4892 2337
rect 4748 2277 4802 2333
rect 4802 2277 4812 2333
rect 4828 2277 4858 2333
rect 4858 2277 4892 2333
rect 4748 2273 4812 2277
rect 4828 2273 4892 2277
rect 4908 2273 4972 2337
rect 4988 2333 5052 2337
rect 5068 2333 5132 2337
rect 4988 2277 5026 2333
rect 5026 2277 5052 2333
rect 5068 2277 5082 2333
rect 5082 2277 5132 2333
rect 4988 2273 5052 2277
rect 5068 2273 5132 2277
rect 5148 2273 5212 2337
rect 5228 2333 5292 2337
rect 5228 2277 5250 2333
rect 5250 2277 5292 2333
rect 5228 2273 5292 2277
rect 5308 2273 5372 2337
rect 5388 2273 5452 2337
rect 5468 2333 5532 2337
rect 5468 2277 5474 2333
rect 5474 2277 5530 2333
rect 5530 2277 5532 2333
rect 5468 2273 5532 2277
rect 5548 2273 5612 2337
rect 5628 2273 5692 2337
rect 5708 2333 5772 2337
rect 5708 2277 5754 2333
rect 5754 2277 5772 2333
rect 5708 2273 5772 2277
rect 5788 2273 5852 2337
rect 5868 2333 5932 2337
rect 5948 2333 6012 2337
rect 5868 2277 5922 2333
rect 5922 2277 5932 2333
rect 5948 2277 5978 2333
rect 5978 2277 6012 2333
rect 5868 2273 5932 2277
rect 5948 2273 6012 2277
rect 6028 2273 6092 2337
rect 6108 2333 6172 2337
rect 6188 2333 6252 2337
rect 6108 2277 6146 2333
rect 6146 2277 6172 2333
rect 6188 2277 6202 2333
rect 6202 2277 6252 2333
rect 6108 2273 6172 2277
rect 6188 2273 6252 2277
rect 6268 2273 6332 2337
rect 6348 2333 6412 2337
rect 6348 2277 6370 2333
rect 6370 2277 6412 2333
rect 6348 2273 6412 2277
rect 6428 2273 6492 2337
rect 6508 2273 6572 2337
rect 6588 2333 6652 2337
rect 6588 2277 6594 2333
rect 6594 2277 6650 2333
rect 6650 2277 6652 2333
rect 6588 2273 6652 2277
rect 6668 2273 6732 2337
rect 6748 2273 6812 2337
rect 6828 2333 6892 2337
rect 6828 2277 6874 2333
rect 6874 2277 6892 2333
rect 6828 2273 6892 2277
rect 6908 2273 6972 2337
rect 6988 2333 7052 2337
rect 7068 2333 7132 2337
rect 6988 2277 7042 2333
rect 7042 2277 7052 2333
rect 7068 2277 7098 2333
rect 7098 2277 7132 2333
rect 6988 2273 7052 2277
rect 7068 2273 7132 2277
rect 7148 2273 7212 2337
rect 7228 2333 7292 2337
rect 7308 2333 7372 2337
rect 7228 2277 7266 2333
rect 7266 2277 7292 2333
rect 7308 2277 7322 2333
rect 7322 2277 7372 2333
rect 7228 2273 7292 2277
rect 7308 2273 7372 2277
rect 7388 2273 7452 2337
rect 7468 2333 7532 2337
rect 7468 2277 7490 2333
rect 7490 2277 7532 2333
rect 7468 2273 7532 2277
rect 7548 2273 7612 2337
rect 7628 2273 7692 2337
rect 7708 2333 7772 2337
rect 7708 2277 7714 2333
rect 7714 2277 7770 2333
rect 7770 2277 7772 2333
rect 7708 2273 7772 2277
rect 7788 2273 7852 2337
rect 7868 2273 7932 2337
rect 7948 2333 8012 2337
rect 7948 2277 7994 2333
rect 7994 2277 8012 2333
rect 7948 2273 8012 2277
rect 8028 2273 8092 2337
rect 8108 2333 8172 2337
rect 8188 2333 8252 2337
rect 8108 2277 8162 2333
rect 8162 2277 8172 2333
rect 8188 2277 8218 2333
rect 8218 2277 8252 2333
rect 8108 2273 8172 2277
rect 8188 2273 8252 2277
rect 8268 2273 8332 2337
rect 8348 2333 8412 2337
rect 8428 2333 8492 2337
rect 8348 2277 8386 2333
rect 8386 2277 8412 2333
rect 8428 2277 8442 2333
rect 8442 2277 8492 2333
rect 8348 2273 8412 2277
rect 8428 2273 8492 2277
rect 8508 2273 8572 2337
rect 8588 2333 8652 2337
rect 8588 2277 8610 2333
rect 8610 2277 8652 2333
rect 8588 2273 8652 2277
rect 8668 2273 8732 2337
rect 8748 2273 8812 2337
rect 8828 2333 8892 2337
rect 8828 2277 8834 2333
rect 8834 2277 8890 2333
rect 8890 2277 8892 2333
rect 8828 2273 8892 2277
rect 8908 2273 8972 2337
rect 8988 2273 9052 2337
rect 9068 2333 9132 2337
rect 9068 2277 9114 2333
rect 9114 2277 9132 2333
rect 9068 2273 9132 2277
rect 9148 2273 9212 2337
rect 9228 2333 9292 2337
rect 9308 2333 9372 2337
rect 9228 2277 9282 2333
rect 9282 2277 9292 2333
rect 9308 2277 9338 2333
rect 9338 2277 9372 2333
rect 9228 2273 9292 2277
rect 9308 2273 9372 2277
rect 9388 2273 9452 2337
rect 9468 2333 9532 2337
rect 9548 2333 9612 2337
rect 9468 2277 9506 2333
rect 9506 2277 9532 2333
rect 9548 2277 9562 2333
rect 9562 2277 9612 2333
rect 9468 2273 9532 2277
rect 9548 2273 9612 2277
rect 9628 2273 9692 2337
rect 9708 2333 9772 2337
rect 9708 2277 9730 2333
rect 9730 2277 9772 2333
rect 9708 2273 9772 2277
rect 9788 2273 9852 2337
rect 9868 2273 9932 2337
rect 9948 2333 10012 2337
rect 9948 2277 9954 2333
rect 9954 2277 10010 2333
rect 10010 2277 10012 2333
rect 9948 2273 10012 2277
rect 10028 2273 10092 2337
rect 10108 2273 10172 2337
rect 10188 2333 10252 2337
rect 10188 2277 10234 2333
rect 10234 2277 10252 2333
rect 10188 2273 10252 2277
rect 10268 2273 10332 2337
rect 10348 2333 10412 2337
rect 10428 2333 10492 2337
rect 10348 2277 10402 2333
rect 10402 2277 10412 2333
rect 10428 2277 10458 2333
rect 10458 2277 10492 2333
rect 10348 2273 10412 2277
rect 10428 2273 10492 2277
rect 10508 2273 10572 2337
rect 10588 2333 10652 2337
rect 10668 2333 10732 2337
rect 10588 2277 10626 2333
rect 10626 2277 10652 2333
rect 10668 2277 10682 2333
rect 10682 2277 10732 2333
rect 10588 2273 10652 2277
rect 10668 2273 10732 2277
rect 10748 2273 10812 2337
rect 10828 2333 10892 2337
rect 10828 2277 10850 2333
rect 10850 2277 10892 2333
rect 10828 2273 10892 2277
rect 10908 2273 10972 2337
rect 10988 2273 11052 2337
rect 28 61 92 65
rect 28 5 42 61
rect 42 5 92 61
rect 28 1 92 5
rect 108 1 172 65
rect 188 1 252 65
rect 268 61 332 65
rect 268 5 322 61
rect 322 5 332 61
rect 268 1 332 5
rect 348 1 412 65
rect 428 61 492 65
rect 508 61 572 65
rect 428 5 490 61
rect 490 5 492 61
rect 508 5 546 61
rect 546 5 572 61
rect 428 1 492 5
rect 508 1 572 5
rect 588 1 652 65
rect 668 61 732 65
rect 748 61 812 65
rect 668 5 714 61
rect 714 5 732 61
rect 748 5 770 61
rect 770 5 812 61
rect 668 1 732 5
rect 748 1 812 5
rect 828 1 892 65
rect 908 61 972 65
rect 988 61 1052 65
rect 908 5 938 61
rect 938 5 972 61
rect 988 5 994 61
rect 994 5 1052 61
rect 908 1 972 5
rect 988 1 1052 5
rect 1068 1 1132 65
rect 1148 61 1212 65
rect 1148 5 1162 61
rect 1162 5 1212 61
rect 1148 1 1212 5
rect 1228 1 1292 65
rect 1308 1 1372 65
rect 1388 61 1452 65
rect 1388 5 1442 61
rect 1442 5 1452 61
rect 1388 1 1452 5
rect 1468 1 1532 65
rect 1548 61 1612 65
rect 1628 61 1692 65
rect 1548 5 1610 61
rect 1610 5 1612 61
rect 1628 5 1666 61
rect 1666 5 1692 61
rect 1548 1 1612 5
rect 1628 1 1692 5
rect 1708 1 1772 65
rect 1788 61 1852 65
rect 1868 61 1932 65
rect 1788 5 1834 61
rect 1834 5 1852 61
rect 1868 5 1890 61
rect 1890 5 1932 61
rect 1788 1 1852 5
rect 1868 1 1932 5
rect 1948 1 2012 65
rect 2028 61 2092 65
rect 2108 61 2172 65
rect 2028 5 2058 61
rect 2058 5 2092 61
rect 2108 5 2114 61
rect 2114 5 2172 61
rect 2028 1 2092 5
rect 2108 1 2172 5
rect 2188 1 2252 65
rect 2268 61 2332 65
rect 2268 5 2282 61
rect 2282 5 2332 61
rect 2268 1 2332 5
rect 2348 1 2412 65
rect 2428 1 2492 65
rect 2508 61 2572 65
rect 2508 5 2562 61
rect 2562 5 2572 61
rect 2508 1 2572 5
rect 2588 1 2652 65
rect 2668 61 2732 65
rect 2748 61 2812 65
rect 2668 5 2730 61
rect 2730 5 2732 61
rect 2748 5 2786 61
rect 2786 5 2812 61
rect 2668 1 2732 5
rect 2748 1 2812 5
rect 2828 1 2892 65
rect 2908 61 2972 65
rect 2988 61 3052 65
rect 2908 5 2954 61
rect 2954 5 2972 61
rect 2988 5 3010 61
rect 3010 5 3052 61
rect 2908 1 2972 5
rect 2988 1 3052 5
rect 3068 1 3132 65
rect 3148 61 3212 65
rect 3228 61 3292 65
rect 3148 5 3178 61
rect 3178 5 3212 61
rect 3228 5 3234 61
rect 3234 5 3292 61
rect 3148 1 3212 5
rect 3228 1 3292 5
rect 3308 1 3372 65
rect 3388 61 3452 65
rect 3388 5 3402 61
rect 3402 5 3452 61
rect 3388 1 3452 5
rect 3468 1 3532 65
rect 3548 1 3612 65
rect 3628 61 3692 65
rect 3628 5 3682 61
rect 3682 5 3692 61
rect 3628 1 3692 5
rect 3708 1 3772 65
rect 3788 61 3852 65
rect 3868 61 3932 65
rect 3788 5 3850 61
rect 3850 5 3852 61
rect 3868 5 3906 61
rect 3906 5 3932 61
rect 3788 1 3852 5
rect 3868 1 3932 5
rect 3948 1 4012 65
rect 4028 61 4092 65
rect 4108 61 4172 65
rect 4028 5 4074 61
rect 4074 5 4092 61
rect 4108 5 4130 61
rect 4130 5 4172 61
rect 4028 1 4092 5
rect 4108 1 4172 5
rect 4188 1 4252 65
rect 4268 61 4332 65
rect 4348 61 4412 65
rect 4268 5 4298 61
rect 4298 5 4332 61
rect 4348 5 4354 61
rect 4354 5 4412 61
rect 4268 1 4332 5
rect 4348 1 4412 5
rect 4428 1 4492 65
rect 4508 61 4572 65
rect 4508 5 4522 61
rect 4522 5 4572 61
rect 4508 1 4572 5
rect 4588 1 4652 65
rect 4668 1 4732 65
rect 4748 61 4812 65
rect 4748 5 4802 61
rect 4802 5 4812 61
rect 4748 1 4812 5
rect 4828 1 4892 65
rect 4908 61 4972 65
rect 4988 61 5052 65
rect 4908 5 4970 61
rect 4970 5 4972 61
rect 4988 5 5026 61
rect 5026 5 5052 61
rect 4908 1 4972 5
rect 4988 1 5052 5
rect 5068 1 5132 65
rect 5148 61 5212 65
rect 5228 61 5292 65
rect 5148 5 5194 61
rect 5194 5 5212 61
rect 5228 5 5250 61
rect 5250 5 5292 61
rect 5148 1 5212 5
rect 5228 1 5292 5
rect 5308 1 5372 65
rect 5388 61 5452 65
rect 5468 61 5532 65
rect 5388 5 5418 61
rect 5418 5 5452 61
rect 5468 5 5474 61
rect 5474 5 5532 61
rect 5388 1 5452 5
rect 5468 1 5532 5
rect 5548 1 5612 65
rect 5628 61 5692 65
rect 5628 5 5642 61
rect 5642 5 5692 61
rect 5628 1 5692 5
rect 5708 1 5772 65
rect 5788 1 5852 65
rect 5868 61 5932 65
rect 5868 5 5922 61
rect 5922 5 5932 61
rect 5868 1 5932 5
rect 5948 1 6012 65
rect 6028 61 6092 65
rect 6108 61 6172 65
rect 6028 5 6090 61
rect 6090 5 6092 61
rect 6108 5 6146 61
rect 6146 5 6172 61
rect 6028 1 6092 5
rect 6108 1 6172 5
rect 6188 1 6252 65
rect 6268 61 6332 65
rect 6348 61 6412 65
rect 6268 5 6314 61
rect 6314 5 6332 61
rect 6348 5 6370 61
rect 6370 5 6412 61
rect 6268 1 6332 5
rect 6348 1 6412 5
rect 6428 1 6492 65
rect 6508 61 6572 65
rect 6588 61 6652 65
rect 6508 5 6538 61
rect 6538 5 6572 61
rect 6588 5 6594 61
rect 6594 5 6652 61
rect 6508 1 6572 5
rect 6588 1 6652 5
rect 6668 1 6732 65
rect 6748 61 6812 65
rect 6748 5 6762 61
rect 6762 5 6812 61
rect 6748 1 6812 5
rect 6828 1 6892 65
rect 6908 1 6972 65
rect 6988 61 7052 65
rect 6988 5 7042 61
rect 7042 5 7052 61
rect 6988 1 7052 5
rect 7068 1 7132 65
rect 7148 61 7212 65
rect 7228 61 7292 65
rect 7148 5 7210 61
rect 7210 5 7212 61
rect 7228 5 7266 61
rect 7266 5 7292 61
rect 7148 1 7212 5
rect 7228 1 7292 5
rect 7308 1 7372 65
rect 7388 61 7452 65
rect 7468 61 7532 65
rect 7388 5 7434 61
rect 7434 5 7452 61
rect 7468 5 7490 61
rect 7490 5 7532 61
rect 7388 1 7452 5
rect 7468 1 7532 5
rect 7548 1 7612 65
rect 7628 61 7692 65
rect 7708 61 7772 65
rect 7628 5 7658 61
rect 7658 5 7692 61
rect 7708 5 7714 61
rect 7714 5 7772 61
rect 7628 1 7692 5
rect 7708 1 7772 5
rect 7788 1 7852 65
rect 7868 61 7932 65
rect 7868 5 7882 61
rect 7882 5 7932 61
rect 7868 1 7932 5
rect 7948 1 8012 65
rect 8028 1 8092 65
rect 8108 61 8172 65
rect 8108 5 8162 61
rect 8162 5 8172 61
rect 8108 1 8172 5
rect 8188 1 8252 65
rect 8268 61 8332 65
rect 8348 61 8412 65
rect 8268 5 8330 61
rect 8330 5 8332 61
rect 8348 5 8386 61
rect 8386 5 8412 61
rect 8268 1 8332 5
rect 8348 1 8412 5
rect 8428 1 8492 65
rect 8508 61 8572 65
rect 8588 61 8652 65
rect 8508 5 8554 61
rect 8554 5 8572 61
rect 8588 5 8610 61
rect 8610 5 8652 61
rect 8508 1 8572 5
rect 8588 1 8652 5
rect 8668 1 8732 65
rect 8748 61 8812 65
rect 8828 61 8892 65
rect 8748 5 8778 61
rect 8778 5 8812 61
rect 8828 5 8834 61
rect 8834 5 8892 61
rect 8748 1 8812 5
rect 8828 1 8892 5
rect 8908 1 8972 65
rect 8988 61 9052 65
rect 8988 5 9002 61
rect 9002 5 9052 61
rect 8988 1 9052 5
rect 9068 1 9132 65
rect 9148 1 9212 65
rect 9228 61 9292 65
rect 9228 5 9282 61
rect 9282 5 9292 61
rect 9228 1 9292 5
rect 9308 1 9372 65
rect 9388 61 9452 65
rect 9468 61 9532 65
rect 9388 5 9450 61
rect 9450 5 9452 61
rect 9468 5 9506 61
rect 9506 5 9532 61
rect 9388 1 9452 5
rect 9468 1 9532 5
rect 9548 1 9612 65
rect 9628 61 9692 65
rect 9708 61 9772 65
rect 9628 5 9674 61
rect 9674 5 9692 61
rect 9708 5 9730 61
rect 9730 5 9772 61
rect 9628 1 9692 5
rect 9708 1 9772 5
rect 9788 1 9852 65
rect 9868 61 9932 65
rect 9948 61 10012 65
rect 9868 5 9898 61
rect 9898 5 9932 61
rect 9948 5 9954 61
rect 9954 5 10012 61
rect 9868 1 9932 5
rect 9948 1 10012 5
rect 10028 1 10092 65
rect 10108 61 10172 65
rect 10108 5 10122 61
rect 10122 5 10172 61
rect 10108 1 10172 5
rect 10188 1 10252 65
rect 10268 1 10332 65
rect 10348 61 10412 65
rect 10348 5 10402 61
rect 10402 5 10412 61
rect 10348 1 10412 5
rect 10428 1 10492 65
rect 10508 61 10572 65
rect 10588 61 10652 65
rect 10508 5 10570 61
rect 10570 5 10572 61
rect 10588 5 10626 61
rect 10626 5 10652 61
rect 10508 1 10572 5
rect 10588 1 10652 5
rect 10668 1 10732 65
rect 10748 61 10812 65
rect 10828 61 10892 65
rect 10748 5 10794 61
rect 10794 5 10812 61
rect 10828 5 10850 61
rect 10850 5 10892 61
rect 10748 1 10812 5
rect 10828 1 10892 5
rect 10908 1 10972 65
rect 10988 61 11052 65
rect 10988 5 11018 61
rect 11018 5 11052 61
rect 10988 1 11052 5
<< metal4 >>
rect 0 2337 11146 2338
rect 0 2273 28 2337
rect 92 2273 108 2337
rect 172 2273 188 2337
rect 252 2273 268 2337
rect 332 2273 348 2337
rect 412 2273 428 2337
rect 492 2273 508 2337
rect 572 2273 588 2337
rect 652 2273 668 2337
rect 732 2273 748 2337
rect 812 2273 828 2337
rect 892 2273 908 2337
rect 972 2273 988 2337
rect 1052 2273 1068 2337
rect 1132 2273 1148 2337
rect 1212 2273 1228 2337
rect 1292 2273 1308 2337
rect 1372 2273 1388 2337
rect 1452 2273 1468 2337
rect 1532 2273 1548 2337
rect 1612 2273 1628 2337
rect 1692 2273 1708 2337
rect 1772 2273 1788 2337
rect 1852 2273 1868 2337
rect 1932 2273 1948 2337
rect 2012 2273 2028 2337
rect 2092 2273 2108 2337
rect 2172 2273 2188 2337
rect 2252 2273 2268 2337
rect 2332 2273 2348 2337
rect 2412 2273 2428 2337
rect 2492 2273 2508 2337
rect 2572 2273 2588 2337
rect 2652 2273 2668 2337
rect 2732 2273 2748 2337
rect 2812 2273 2828 2337
rect 2892 2273 2908 2337
rect 2972 2273 2988 2337
rect 3052 2273 3068 2337
rect 3132 2273 3148 2337
rect 3212 2273 3228 2337
rect 3292 2273 3308 2337
rect 3372 2273 3388 2337
rect 3452 2273 3468 2337
rect 3532 2273 3548 2337
rect 3612 2273 3628 2337
rect 3692 2273 3708 2337
rect 3772 2273 3788 2337
rect 3852 2273 3868 2337
rect 3932 2273 3948 2337
rect 4012 2273 4028 2337
rect 4092 2273 4108 2337
rect 4172 2273 4188 2337
rect 4252 2273 4268 2337
rect 4332 2273 4348 2337
rect 4412 2273 4428 2337
rect 4492 2273 4508 2337
rect 4572 2273 4588 2337
rect 4652 2273 4668 2337
rect 4732 2273 4748 2337
rect 4812 2273 4828 2337
rect 4892 2273 4908 2337
rect 4972 2273 4988 2337
rect 5052 2273 5068 2337
rect 5132 2273 5148 2337
rect 5212 2273 5228 2337
rect 5292 2273 5308 2337
rect 5372 2273 5388 2337
rect 5452 2273 5468 2337
rect 5532 2273 5548 2337
rect 5612 2273 5628 2337
rect 5692 2273 5708 2337
rect 5772 2273 5788 2337
rect 5852 2273 5868 2337
rect 5932 2273 5948 2337
rect 6012 2273 6028 2337
rect 6092 2273 6108 2337
rect 6172 2273 6188 2337
rect 6252 2273 6268 2337
rect 6332 2273 6348 2337
rect 6412 2273 6428 2337
rect 6492 2273 6508 2337
rect 6572 2273 6588 2337
rect 6652 2273 6668 2337
rect 6732 2273 6748 2337
rect 6812 2273 6828 2337
rect 6892 2273 6908 2337
rect 6972 2273 6988 2337
rect 7052 2273 7068 2337
rect 7132 2273 7148 2337
rect 7212 2273 7228 2337
rect 7292 2273 7308 2337
rect 7372 2273 7388 2337
rect 7452 2273 7468 2337
rect 7532 2273 7548 2337
rect 7612 2273 7628 2337
rect 7692 2273 7708 2337
rect 7772 2273 7788 2337
rect 7852 2273 7868 2337
rect 7932 2273 7948 2337
rect 8012 2273 8028 2337
rect 8092 2273 8108 2337
rect 8172 2273 8188 2337
rect 8252 2273 8268 2337
rect 8332 2273 8348 2337
rect 8412 2273 8428 2337
rect 8492 2273 8508 2337
rect 8572 2273 8588 2337
rect 8652 2273 8668 2337
rect 8732 2273 8748 2337
rect 8812 2273 8828 2337
rect 8892 2273 8908 2337
rect 8972 2273 8988 2337
rect 9052 2273 9068 2337
rect 9132 2273 9148 2337
rect 9212 2273 9228 2337
rect 9292 2273 9308 2337
rect 9372 2273 9388 2337
rect 9452 2273 9468 2337
rect 9532 2273 9548 2337
rect 9612 2273 9628 2337
rect 9692 2273 9708 2337
rect 9772 2273 9788 2337
rect 9852 2273 9868 2337
rect 9932 2273 9948 2337
rect 10012 2273 10028 2337
rect 10092 2273 10108 2337
rect 10172 2273 10188 2337
rect 10252 2273 10268 2337
rect 10332 2273 10348 2337
rect 10412 2273 10428 2337
rect 10492 2273 10508 2337
rect 10572 2273 10588 2337
rect 10652 2273 10668 2337
rect 10732 2273 10748 2337
rect 10812 2273 10828 2337
rect 10892 2273 10908 2337
rect 10972 2273 10988 2337
rect 11052 2273 11146 2337
rect 0 2272 11146 2273
rect 120 2234 420 2272
rect 0 66 60 2212
rect 120 1998 152 2234
rect 388 1998 420 2234
rect 120 126 180 1998
rect 240 340 300 1938
rect 360 400 420 1998
rect 480 340 540 2212
rect 240 104 272 340
rect 508 104 540 340
rect 600 126 660 2272
rect 240 66 540 104
rect 720 66 780 2212
rect 840 126 900 2272
rect 960 66 1020 2212
rect 1080 126 1140 2272
rect 1200 66 1260 2212
rect 1320 126 1380 2272
rect 1560 2234 1860 2272
rect 1440 66 1500 2212
rect 1560 1998 1592 2234
rect 1828 1998 1860 2234
rect 1560 126 1620 1998
rect 1680 340 1740 1938
rect 1800 400 1860 1998
rect 1920 340 1980 2212
rect 1680 104 1712 340
rect 1948 104 1980 340
rect 2040 126 2100 2272
rect 1680 66 1980 104
rect 2160 66 2220 2212
rect 2280 126 2340 2272
rect 2400 66 2460 2212
rect 2520 126 2580 2272
rect 2640 66 2700 2212
rect 2760 126 2820 2272
rect 3000 2234 3300 2272
rect 2880 66 2940 2212
rect 3000 1998 3032 2234
rect 3268 1998 3300 2234
rect 3000 126 3060 1998
rect 3120 340 3180 1938
rect 3240 400 3300 1998
rect 3360 340 3420 2212
rect 3120 104 3152 340
rect 3388 104 3420 340
rect 3480 126 3540 2272
rect 3120 66 3420 104
rect 3600 66 3660 2212
rect 3720 126 3780 2272
rect 3840 66 3900 2212
rect 3960 126 4020 2272
rect 4080 66 4140 2212
rect 4200 126 4260 2272
rect 4440 2234 4740 2272
rect 4320 66 4380 2212
rect 4440 1998 4472 2234
rect 4708 1998 4740 2234
rect 4440 126 4500 1998
rect 4560 340 4620 1938
rect 4680 400 4740 1998
rect 4800 340 4860 2212
rect 4560 104 4592 340
rect 4828 104 4860 340
rect 4920 126 4980 2272
rect 4560 66 4860 104
rect 5040 66 5100 2212
rect 5160 126 5220 2272
rect 5280 66 5340 2212
rect 5400 126 5460 2272
rect 5520 66 5580 2212
rect 5640 126 5700 2272
rect 5880 2234 6180 2272
rect 5760 66 5820 2212
rect 5880 1998 5912 2234
rect 6148 1998 6180 2234
rect 5880 126 5940 1998
rect 6000 340 6060 1938
rect 6120 400 6180 1998
rect 6240 340 6300 2212
rect 6000 104 6032 340
rect 6268 104 6300 340
rect 6360 126 6420 2272
rect 6000 66 6300 104
rect 6480 66 6540 2212
rect 6600 126 6660 2272
rect 6720 66 6780 2212
rect 6840 126 6900 2272
rect 6960 66 7020 2212
rect 7080 126 7140 2272
rect 7320 2234 7620 2272
rect 7200 66 7260 2212
rect 7320 1998 7352 2234
rect 7588 1998 7620 2234
rect 7320 126 7380 1998
rect 7440 340 7500 1938
rect 7560 400 7620 1998
rect 7680 340 7740 2212
rect 7440 104 7472 340
rect 7708 104 7740 340
rect 7800 126 7860 2272
rect 7440 66 7740 104
rect 7920 66 7980 2212
rect 8040 126 8100 2272
rect 8160 66 8220 2212
rect 8280 126 8340 2272
rect 8400 66 8460 2212
rect 8520 126 8580 2272
rect 8760 2234 9060 2272
rect 8640 66 8700 2212
rect 8760 1998 8792 2234
rect 9028 1998 9060 2234
rect 8760 126 8820 1998
rect 8880 340 8940 1938
rect 9000 400 9060 1998
rect 9120 340 9180 2212
rect 8880 104 8912 340
rect 9148 104 9180 340
rect 9240 126 9300 2272
rect 8880 66 9180 104
rect 9360 66 9420 2212
rect 9480 126 9540 2272
rect 9600 66 9660 2212
rect 9720 126 9780 2272
rect 9840 66 9900 2212
rect 9960 126 10020 2272
rect 10200 2234 10500 2272
rect 10080 66 10140 2212
rect 10200 1998 10232 2234
rect 10468 1998 10500 2234
rect 10200 126 10260 1998
rect 10320 340 10380 1938
rect 10440 400 10500 1998
rect 10560 340 10620 2212
rect 10320 104 10352 340
rect 10588 104 10620 340
rect 10680 126 10740 2272
rect 10320 66 10620 104
rect 10800 66 10860 2212
rect 10920 126 10980 2272
rect 11040 66 11146 2212
rect 0 65 11146 66
rect 0 1 28 65
rect 92 1 108 65
rect 172 1 188 65
rect 252 1 268 65
rect 332 1 348 65
rect 412 1 428 65
rect 492 1 508 65
rect 572 1 588 65
rect 652 1 668 65
rect 732 1 748 65
rect 812 1 828 65
rect 892 1 908 65
rect 972 1 988 65
rect 1052 1 1068 65
rect 1132 1 1148 65
rect 1212 1 1228 65
rect 1292 1 1308 65
rect 1372 1 1388 65
rect 1452 1 1468 65
rect 1532 1 1548 65
rect 1612 1 1628 65
rect 1692 1 1708 65
rect 1772 1 1788 65
rect 1852 1 1868 65
rect 1932 1 1948 65
rect 2012 1 2028 65
rect 2092 1 2108 65
rect 2172 1 2188 65
rect 2252 1 2268 65
rect 2332 1 2348 65
rect 2412 1 2428 65
rect 2492 1 2508 65
rect 2572 1 2588 65
rect 2652 1 2668 65
rect 2732 1 2748 65
rect 2812 1 2828 65
rect 2892 1 2908 65
rect 2972 1 2988 65
rect 3052 1 3068 65
rect 3132 1 3148 65
rect 3212 1 3228 65
rect 3292 1 3308 65
rect 3372 1 3388 65
rect 3452 1 3468 65
rect 3532 1 3548 65
rect 3612 1 3628 65
rect 3692 1 3708 65
rect 3772 1 3788 65
rect 3852 1 3868 65
rect 3932 1 3948 65
rect 4012 1 4028 65
rect 4092 1 4108 65
rect 4172 1 4188 65
rect 4252 1 4268 65
rect 4332 1 4348 65
rect 4412 1 4428 65
rect 4492 1 4508 65
rect 4572 1 4588 65
rect 4652 1 4668 65
rect 4732 1 4748 65
rect 4812 1 4828 65
rect 4892 1 4908 65
rect 4972 1 4988 65
rect 5052 1 5068 65
rect 5132 1 5148 65
rect 5212 1 5228 65
rect 5292 1 5308 65
rect 5372 1 5388 65
rect 5452 1 5468 65
rect 5532 1 5548 65
rect 5612 1 5628 65
rect 5692 1 5708 65
rect 5772 1 5788 65
rect 5852 1 5868 65
rect 5932 1 5948 65
rect 6012 1 6028 65
rect 6092 1 6108 65
rect 6172 1 6188 65
rect 6252 1 6268 65
rect 6332 1 6348 65
rect 6412 1 6428 65
rect 6492 1 6508 65
rect 6572 1 6588 65
rect 6652 1 6668 65
rect 6732 1 6748 65
rect 6812 1 6828 65
rect 6892 1 6908 65
rect 6972 1 6988 65
rect 7052 1 7068 65
rect 7132 1 7148 65
rect 7212 1 7228 65
rect 7292 1 7308 65
rect 7372 1 7388 65
rect 7452 1 7468 65
rect 7532 1 7548 65
rect 7612 1 7628 65
rect 7692 1 7708 65
rect 7772 1 7788 65
rect 7852 1 7868 65
rect 7932 1 7948 65
rect 8012 1 8028 65
rect 8092 1 8108 65
rect 8172 1 8188 65
rect 8252 1 8268 65
rect 8332 1 8348 65
rect 8412 1 8428 65
rect 8492 1 8508 65
rect 8572 1 8588 65
rect 8652 1 8668 65
rect 8732 1 8748 65
rect 8812 1 8828 65
rect 8892 1 8908 65
rect 8972 1 8988 65
rect 9052 1 9068 65
rect 9132 1 9148 65
rect 9212 1 9228 65
rect 9292 1 9308 65
rect 9372 1 9388 65
rect 9452 1 9468 65
rect 9532 1 9548 65
rect 9612 1 9628 65
rect 9692 1 9708 65
rect 9772 1 9788 65
rect 9852 1 9868 65
rect 9932 1 9948 65
rect 10012 1 10028 65
rect 10092 1 10108 65
rect 10172 1 10188 65
rect 10252 1 10268 65
rect 10332 1 10348 65
rect 10412 1 10428 65
rect 10492 1 10508 65
rect 10572 1 10588 65
rect 10652 1 10668 65
rect 10732 1 10748 65
rect 10812 1 10828 65
rect 10892 1 10908 65
rect 10972 1 10988 65
rect 11052 1 11146 65
rect 0 0 11146 1
<< via4 >>
rect 152 1998 388 2234
rect 272 104 508 340
rect 1592 1998 1828 2234
rect 1712 104 1948 340
rect 3032 1998 3268 2234
rect 3152 104 3388 340
rect 4472 1998 4708 2234
rect 4592 104 4828 340
rect 5912 1998 6148 2234
rect 6032 104 6268 340
rect 7352 1998 7588 2234
rect 7472 104 7708 340
rect 8792 1998 9028 2234
rect 8912 104 9148 340
rect 10232 1998 10468 2234
rect 10352 104 10588 340
<< metal5 >>
rect 0 2234 10986 2258
rect 0 1998 152 2234
rect 388 1998 1592 2234
rect 1828 1998 3032 2234
rect 3268 1998 4472 2234
rect 4708 1998 5912 2234
rect 6148 1998 7352 2234
rect 7588 1998 8792 2234
rect 9028 1998 10232 2234
rect 10468 1998 10986 2234
rect 0 1938 10986 1998
rect 0 720 320 1938
rect 640 400 960 1618
rect 1280 720 1600 1938
rect 1920 400 2240 1618
rect 2560 720 2880 1938
rect 3200 400 3520 1618
rect 3840 720 4160 1938
rect 4480 400 4800 1618
rect 5120 720 5440 1938
rect 5760 400 6080 1618
rect 6400 720 6720 1938
rect 7040 400 7360 1618
rect 7680 720 8000 1938
rect 8320 400 8640 1618
rect 8960 720 9280 1938
rect 9600 400 9920 1618
rect 10240 720 10986 1938
rect 0 340 10986 400
rect 0 104 272 340
rect 508 104 1712 340
rect 1948 104 3152 340
rect 3388 104 4592 340
rect 4828 104 6032 340
rect 6268 104 7472 340
rect 7708 104 8912 340
rect 9148 104 10352 340
rect 10588 104 10986 340
rect 0 80 10986 104
<< properties >>
string GDS_END 2155188
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 1999152
<< end >>
