magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 827 203
rect 30 -17 64 21
<< locali >>
rect 103 59 169 485
rect 299 199 342 265
rect 379 121 433 265
rect 488 199 535 265
rect 579 199 647 265
rect 739 199 801 265
rect 488 121 524 199
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 299 69 527
rect 18 17 69 177
rect 232 367 276 527
rect 318 401 368 493
rect 425 451 491 527
rect 543 401 605 493
rect 318 367 605 401
rect 759 333 793 493
rect 203 299 793 333
rect 203 165 237 299
rect 203 131 339 165
rect 203 17 269 93
rect 305 85 339 131
rect 558 131 793 165
rect 558 85 592 131
rect 305 51 592 85
rect 644 17 710 97
rect 759 51 793 131
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 488 121 524 199 6 A1
port 1 nsew signal input
rlabel locali s 488 199 535 265 6 A1
port 1 nsew signal input
rlabel locali s 379 121 433 265 6 A2
port 2 nsew signal input
rlabel locali s 299 199 342 265 6 A3
port 3 nsew signal input
rlabel locali s 579 199 647 265 6 B1
port 4 nsew signal input
rlabel locali s 739 199 801 265 6 C1
port 5 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 827 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 103 59 169 485 6 X
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3708814
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3701494
<< end >>
