magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< locali >>
rect 0 527 736 561
rect 0 -17 736 17
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 0 -17 736 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 0 527 736 561 6 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 496 736 592 6 VPWR
port 2 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE SPACER
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3952840
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3950588
<< end >>
