magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -66 377 2466 897
<< pwell >>
rect 2134 289 2396 317
rect 4 223 426 237
rect 1153 223 1435 289
rect 1862 223 2396 289
rect 4 43 2396 223
rect -26 -43 2426 43
<< mvnmos >>
rect 87 127 187 211
rect 243 127 343 211
rect 540 113 640 197
rect 720 113 820 197
rect 915 113 1015 197
rect 1057 113 1157 197
rect 1252 113 1352 263
rect 1431 113 1531 197
rect 1587 113 1687 197
rect 1729 113 1829 197
rect 1941 113 2041 263
rect 2217 141 2317 291
<< mvpmos >>
rect 83 559 183 709
rect 239 559 339 709
rect 505 563 605 647
rect 680 574 780 658
rect 882 543 982 627
rect 1024 543 1124 627
rect 1199 543 1299 743
rect 1355 543 1455 743
rect 1631 543 1731 627
rect 1773 543 1873 627
rect 1948 543 2048 743
rect 2217 443 2317 743
<< mvndiff >>
rect 30 186 87 211
rect 30 152 42 186
rect 76 152 87 186
rect 30 127 87 152
rect 187 186 243 211
rect 187 152 198 186
rect 232 152 243 186
rect 187 127 243 152
rect 343 186 400 211
rect 1179 197 1252 263
rect 343 152 354 186
rect 388 152 400 186
rect 343 127 400 152
rect 483 172 540 197
rect 483 138 495 172
rect 529 138 540 172
rect 483 113 540 138
rect 640 173 720 197
rect 640 139 675 173
rect 709 139 720 173
rect 640 113 720 139
rect 820 173 915 197
rect 820 139 859 173
rect 893 139 915 173
rect 820 113 915 139
rect 1015 113 1057 197
rect 1157 177 1252 197
rect 1157 143 1191 177
rect 1225 143 1252 177
rect 1157 113 1252 143
rect 1352 255 1409 263
rect 1352 221 1363 255
rect 1397 221 1409 255
rect 1352 197 1409 221
rect 2160 283 2217 291
rect 1888 249 1941 263
rect 1888 215 1896 249
rect 1930 215 1941 249
rect 1888 197 1941 215
rect 1352 157 1431 197
rect 1352 123 1363 157
rect 1397 123 1431 157
rect 1352 113 1431 123
rect 1531 172 1587 197
rect 1531 138 1542 172
rect 1576 138 1587 172
rect 1531 113 1587 138
rect 1687 113 1729 197
rect 1829 159 1941 197
rect 1829 125 1896 159
rect 1930 125 1941 159
rect 1829 113 1941 125
rect 2041 255 2098 263
rect 2041 221 2052 255
rect 2086 221 2098 255
rect 2041 155 2098 221
rect 2041 121 2052 155
rect 2086 121 2098 155
rect 2160 249 2172 283
rect 2206 249 2217 283
rect 2160 183 2217 249
rect 2160 149 2172 183
rect 2206 149 2217 183
rect 2160 141 2217 149
rect 2317 279 2370 291
rect 2317 245 2328 279
rect 2362 245 2370 279
rect 2317 187 2370 245
rect 2317 153 2328 187
rect 2362 153 2370 187
rect 2317 141 2370 153
rect 2041 113 2098 121
<< mvpdiff >>
rect 1146 731 1199 743
rect 30 697 83 709
rect 30 663 38 697
rect 72 663 83 697
rect 30 605 83 663
rect 30 571 38 605
rect 72 571 83 605
rect 30 559 83 571
rect 183 701 239 709
rect 183 667 194 701
rect 228 667 239 701
rect 183 601 239 667
rect 183 567 194 601
rect 228 567 239 601
rect 183 559 239 567
rect 339 697 392 709
rect 339 663 350 697
rect 384 663 392 697
rect 1146 697 1154 731
rect 1188 697 1199 731
rect 339 605 392 663
rect 630 647 680 658
rect 339 571 350 605
rect 384 571 392 605
rect 339 559 392 571
rect 452 622 505 647
rect 452 588 460 622
rect 494 588 505 622
rect 452 563 505 588
rect 605 617 680 647
rect 605 583 616 617
rect 650 583 680 617
rect 605 574 680 583
rect 780 627 860 658
rect 1146 627 1199 697
rect 780 588 882 627
rect 780 574 827 588
rect 605 563 658 574
rect 802 554 827 574
rect 861 554 882 588
rect 802 543 882 554
rect 982 543 1024 627
rect 1124 543 1199 627
rect 1299 588 1355 743
rect 1299 554 1310 588
rect 1344 554 1355 588
rect 1299 543 1355 554
rect 1455 731 1609 743
rect 1455 697 1567 731
rect 1601 697 1609 731
rect 1455 660 1609 697
rect 1455 626 1567 660
rect 1601 627 1609 660
rect 1895 731 1948 743
rect 1895 697 1903 731
rect 1937 697 1948 731
rect 1895 660 1948 697
rect 1895 627 1903 660
rect 1601 626 1631 627
rect 1455 589 1631 626
rect 1455 555 1567 589
rect 1601 555 1631 589
rect 1455 543 1631 555
rect 1731 543 1773 627
rect 1873 626 1903 627
rect 1937 626 1948 660
rect 1873 589 1948 626
rect 1873 555 1903 589
rect 1937 555 1948 589
rect 1873 543 1948 555
rect 2048 731 2101 743
rect 2048 697 2059 731
rect 2093 697 2101 731
rect 2048 660 2101 697
rect 2048 626 2059 660
rect 2093 626 2101 660
rect 2048 589 2101 626
rect 2048 555 2059 589
rect 2093 555 2101 589
rect 2048 543 2101 555
rect 2164 731 2217 743
rect 2164 697 2172 731
rect 2206 697 2217 731
rect 2164 651 2217 697
rect 2164 617 2172 651
rect 2206 617 2217 651
rect 2164 569 2217 617
rect 2164 535 2172 569
rect 2206 535 2217 569
rect 2164 489 2217 535
rect 2164 455 2172 489
rect 2206 455 2217 489
rect 2164 443 2217 455
rect 2317 731 2370 743
rect 2317 697 2328 731
rect 2362 697 2370 731
rect 2317 651 2370 697
rect 2317 617 2328 651
rect 2362 617 2370 651
rect 2317 569 2370 617
rect 2317 535 2328 569
rect 2362 535 2370 569
rect 2317 489 2370 535
rect 2317 455 2328 489
rect 2362 455 2370 489
rect 2317 443 2370 455
<< mvndiffc >>
rect 42 152 76 186
rect 198 152 232 186
rect 354 152 388 186
rect 495 138 529 172
rect 675 139 709 173
rect 859 139 893 173
rect 1191 143 1225 177
rect 1363 221 1397 255
rect 1896 215 1930 249
rect 1363 123 1397 157
rect 1542 138 1576 172
rect 1896 125 1930 159
rect 2052 221 2086 255
rect 2052 121 2086 155
rect 2172 249 2206 283
rect 2172 149 2206 183
rect 2328 245 2362 279
rect 2328 153 2362 187
<< mvpdiffc >>
rect 38 663 72 697
rect 38 571 72 605
rect 194 667 228 701
rect 194 567 228 601
rect 350 663 384 697
rect 1154 697 1188 731
rect 350 571 384 605
rect 460 588 494 622
rect 616 583 650 617
rect 827 554 861 588
rect 1310 554 1344 588
rect 1567 697 1601 731
rect 1567 626 1601 660
rect 1903 697 1937 731
rect 1567 555 1601 589
rect 1903 626 1937 660
rect 1903 555 1937 589
rect 2059 697 2093 731
rect 2059 626 2093 660
rect 2059 555 2093 589
rect 2172 697 2206 731
rect 2172 617 2206 651
rect 2172 535 2206 569
rect 2172 455 2206 489
rect 2328 697 2362 731
rect 2328 617 2362 651
rect 2328 535 2362 569
rect 2328 455 2362 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2400 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
<< poly >>
rect 1199 743 1299 769
rect 1355 743 1455 769
rect 1948 743 2048 769
rect 2217 743 2317 769
rect 83 709 183 735
rect 239 709 339 735
rect 505 647 605 673
rect 680 658 780 684
rect 882 627 982 653
rect 1024 627 1124 653
rect 83 533 183 559
rect 239 533 339 559
rect 505 537 605 563
rect 83 499 187 533
rect 83 465 124 499
rect 158 465 187 499
rect 83 431 187 465
rect 83 397 124 431
rect 158 397 187 431
rect 83 233 187 397
rect 229 449 339 533
rect 229 429 343 449
rect 229 395 249 429
rect 283 395 343 429
rect 229 361 343 395
rect 229 327 249 361
rect 283 327 343 361
rect 229 237 343 327
rect 424 437 605 537
rect 680 526 780 574
rect 1631 627 1731 653
rect 1773 627 1873 653
rect 680 492 718 526
rect 752 492 780 526
rect 882 517 982 543
rect 680 448 780 492
rect 822 495 982 517
rect 822 461 928 495
rect 962 461 982 495
rect 424 368 540 437
rect 822 427 982 461
rect 822 393 928 427
rect 962 393 982 427
rect 822 379 982 393
rect 682 373 982 379
rect 1024 517 1124 543
rect 1024 425 1157 517
rect 1024 391 1103 425
rect 1137 391 1157 425
rect 424 348 640 368
rect 424 314 444 348
rect 478 314 640 348
rect 424 268 640 314
rect 87 211 187 233
rect 243 211 343 237
rect 540 197 640 268
rect 682 359 867 373
rect 1024 371 1157 391
rect 682 325 702 359
rect 736 325 867 359
rect 682 291 867 325
rect 682 257 702 291
rect 736 257 867 291
rect 682 223 867 257
rect 915 269 1015 319
rect 915 235 961 269
rect 995 235 1015 269
rect 720 197 820 223
rect 915 197 1015 235
rect 1057 197 1157 371
rect 1199 382 1299 543
rect 1355 521 1455 543
rect 1631 521 1731 543
rect 1341 495 1500 521
rect 1341 461 1357 495
rect 1391 461 1500 495
rect 1341 424 1500 461
rect 1580 495 1731 521
rect 1580 461 1600 495
rect 1634 461 1731 495
rect 1580 445 1731 461
rect 1400 403 1500 424
rect 1773 403 1873 543
rect 1948 493 2048 543
rect 1199 339 1352 382
rect 1199 305 1219 339
rect 1253 305 1352 339
rect 1400 335 1681 403
rect 1729 387 1873 403
rect 1729 353 1816 387
rect 1850 353 1873 387
rect 1199 285 1352 305
rect 1252 263 1352 285
rect 1431 273 1531 293
rect 87 101 187 127
rect 243 101 343 127
rect 1431 239 1472 273
rect 1506 239 1531 273
rect 1431 197 1531 239
rect 1581 223 1687 335
rect 1587 197 1687 223
rect 1729 319 1873 353
rect 1937 473 2048 493
rect 1937 439 1957 473
rect 1991 439 2048 473
rect 1937 405 2048 439
rect 2217 417 2317 443
rect 1937 371 1957 405
rect 1991 371 2048 405
rect 1937 351 2048 371
rect 1729 285 1816 319
rect 1850 285 1873 319
rect 1729 265 1873 285
rect 1941 289 2048 351
rect 2090 385 2317 417
rect 2090 351 2106 385
rect 2140 351 2174 385
rect 2208 351 2242 385
rect 2276 351 2317 385
rect 2090 317 2317 351
rect 2217 291 2317 317
rect 1729 197 1829 265
rect 1941 263 2041 289
rect 2217 115 2317 141
rect 540 87 640 113
rect 720 87 820 113
rect 915 87 1015 113
rect 1057 87 1157 113
rect 1252 87 1352 113
rect 1431 87 1531 113
rect 1587 87 1687 113
rect 1729 87 1829 113
rect 1941 87 2041 113
<< polycont >>
rect 124 465 158 499
rect 124 397 158 431
rect 249 395 283 429
rect 249 327 283 361
rect 718 492 752 526
rect 928 461 962 495
rect 928 393 962 427
rect 1103 391 1137 425
rect 444 314 478 348
rect 702 325 736 359
rect 702 257 736 291
rect 961 235 995 269
rect 1357 461 1391 495
rect 1600 461 1634 495
rect 1219 305 1253 339
rect 1816 353 1850 387
rect 1472 239 1506 273
rect 1957 439 1991 473
rect 1957 371 1991 405
rect 1816 285 1850 319
rect 2106 351 2140 385
rect 2174 351 2208 385
rect 2242 351 2276 385
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2400 831
rect 108 735 298 741
rect 22 697 72 713
rect 22 663 38 697
rect 22 605 72 663
rect 22 571 38 605
rect 22 345 72 571
rect 108 701 114 735
rect 148 701 186 735
rect 220 701 258 735
rect 292 701 298 735
rect 444 735 494 741
rect 108 667 194 701
rect 228 667 298 701
rect 108 601 298 667
rect 108 567 194 601
rect 228 567 298 601
rect 108 551 298 567
rect 334 697 400 713
rect 334 663 350 697
rect 384 663 400 697
rect 334 605 400 663
rect 334 571 350 605
rect 384 571 400 605
rect 334 523 400 571
rect 444 701 450 735
rect 484 701 494 735
rect 444 622 494 701
rect 1014 737 1204 747
rect 1014 703 1020 737
rect 1054 703 1092 737
rect 1126 731 1164 737
rect 1126 703 1154 731
rect 1198 703 1204 737
rect 1014 697 1154 703
rect 1188 697 1204 703
rect 1567 731 1617 747
rect 1601 697 1617 731
rect 444 588 460 622
rect 444 559 494 588
rect 530 661 736 695
rect 530 523 564 661
rect 702 627 1531 661
rect 108 499 174 515
rect 108 465 124 499
rect 158 465 174 499
rect 334 489 564 523
rect 600 617 666 625
rect 600 583 616 617
rect 650 583 666 617
rect 108 431 174 465
rect 600 456 666 583
rect 702 526 768 627
rect 811 588 877 591
rect 811 554 827 588
rect 861 554 877 588
rect 811 535 877 554
rect 1294 588 1461 591
rect 1294 554 1310 588
rect 1344 554 1461 588
rect 1294 551 1461 554
rect 702 492 718 526
rect 752 492 768 526
rect 108 397 124 431
rect 158 397 174 431
rect 108 381 174 397
rect 233 429 564 445
rect 233 395 249 429
rect 283 395 564 429
rect 600 422 807 456
rect 233 386 564 395
rect 233 361 283 386
rect 233 345 249 361
rect 22 327 249 345
rect 530 359 737 386
rect 530 352 702 359
rect 22 311 283 327
rect 319 348 494 350
rect 319 314 444 348
rect 478 314 494 348
rect 319 311 494 314
rect 686 325 702 352
rect 736 325 737 359
rect 22 186 76 311
rect 686 291 737 325
rect 338 241 623 275
rect 686 257 702 291
rect 736 257 737 291
rect 686 241 737 257
rect 22 152 42 186
rect 22 119 76 152
rect 112 186 302 219
rect 112 152 198 186
rect 232 152 302 186
rect 112 113 302 152
rect 338 186 404 241
rect 338 152 354 186
rect 388 152 404 186
rect 338 119 404 152
rect 440 172 553 205
rect 440 138 495 172
rect 529 138 553 172
rect 112 79 118 113
rect 152 79 190 113
rect 224 79 262 113
rect 296 79 302 113
rect 112 73 302 79
rect 440 113 553 138
rect 440 79 443 113
rect 477 79 515 113
rect 549 79 553 113
rect 440 73 553 79
rect 589 87 623 241
rect 773 205 807 422
rect 659 173 807 205
rect 659 139 675 173
rect 709 139 807 173
rect 659 123 807 139
rect 843 339 877 535
rect 913 495 1391 511
rect 913 461 928 495
rect 962 477 1357 495
rect 962 461 978 477
rect 913 427 978 461
rect 1341 461 1357 477
rect 1341 445 1391 461
rect 913 393 928 427
rect 962 393 978 427
rect 913 377 978 393
rect 1087 425 1153 441
rect 1087 391 1103 425
rect 1137 409 1153 425
rect 1427 409 1461 551
rect 1137 391 1461 409
rect 1087 375 1461 391
rect 1497 503 1531 627
rect 1567 660 1617 697
rect 1601 626 1617 660
rect 1567 589 1617 626
rect 1601 573 1617 589
rect 1763 735 1953 747
rect 1763 701 1769 735
rect 1803 701 1841 735
rect 1875 731 1913 735
rect 1875 701 1903 731
rect 1947 701 1953 735
rect 1763 697 1903 701
rect 1937 697 1953 701
rect 1763 660 1953 697
rect 1763 626 1903 660
rect 1937 626 1953 660
rect 1763 589 1953 626
rect 1601 555 1720 573
rect 1567 539 1720 555
rect 1763 555 1903 589
rect 1937 555 1953 589
rect 1763 539 1953 555
rect 2043 731 2109 747
rect 2043 697 2059 731
rect 2093 697 2109 731
rect 2043 660 2109 697
rect 2043 626 2059 660
rect 2093 626 2109 660
rect 2043 589 2109 626
rect 2043 555 2059 589
rect 2093 555 2109 589
rect 1497 495 1650 503
rect 1497 461 1600 495
rect 1634 461 1650 495
rect 1497 445 1650 461
rect 1686 489 1720 539
rect 1686 473 2007 489
rect 1686 455 1957 473
rect 843 305 1219 339
rect 1253 305 1269 339
rect 843 173 909 305
rect 843 139 859 173
rect 893 139 909 173
rect 843 123 909 139
rect 945 235 961 269
rect 995 235 1311 269
rect 945 87 1011 235
rect 589 53 1011 87
rect 1051 177 1241 199
rect 1051 143 1191 177
rect 1225 143 1241 177
rect 1051 113 1241 143
rect 1051 79 1057 113
rect 1091 79 1129 113
rect 1163 79 1201 113
rect 1235 79 1241 113
rect 1051 73 1241 79
rect 1277 87 1311 235
rect 1347 255 1413 375
rect 1497 289 1531 445
rect 1347 221 1363 255
rect 1397 221 1413 255
rect 1347 157 1413 221
rect 1347 123 1363 157
rect 1397 123 1413 157
rect 1456 273 1531 289
rect 1456 239 1472 273
rect 1506 239 1531 273
rect 1456 225 1531 239
rect 1456 87 1490 225
rect 1686 205 1720 455
rect 1941 439 1957 455
rect 1991 439 2007 473
rect 1941 405 2007 439
rect 1800 387 1866 403
rect 1800 353 1816 387
rect 1850 353 1866 387
rect 1941 371 1957 405
rect 1991 371 2007 405
rect 1941 355 2007 371
rect 2043 401 2109 555
rect 2145 735 2263 747
rect 2145 701 2151 735
rect 2185 731 2223 735
rect 2206 701 2223 731
rect 2257 701 2263 735
rect 2145 697 2172 701
rect 2206 697 2263 701
rect 2145 651 2263 697
rect 2145 617 2172 651
rect 2206 617 2263 651
rect 2145 569 2263 617
rect 2145 535 2172 569
rect 2206 535 2263 569
rect 2145 489 2263 535
rect 2145 455 2172 489
rect 2206 455 2263 489
rect 2145 439 2263 455
rect 2312 731 2378 747
rect 2312 697 2328 731
rect 2362 697 2378 731
rect 2312 651 2378 697
rect 2312 617 2328 651
rect 2362 617 2378 651
rect 2312 569 2378 617
rect 2312 535 2328 569
rect 2362 535 2378 569
rect 2312 489 2378 535
rect 2312 455 2328 489
rect 2362 455 2378 489
rect 2312 437 2378 455
rect 2043 385 2292 401
rect 1800 319 1866 353
rect 2043 351 2106 385
rect 2140 351 2174 385
rect 2208 351 2242 385
rect 2276 351 2292 385
rect 2043 335 2292 351
rect 2043 319 2102 335
rect 1800 285 1816 319
rect 1850 285 2102 319
rect 2036 255 2102 285
rect 1567 189 1720 205
rect 1526 172 1720 189
rect 1526 138 1542 172
rect 1576 171 1720 172
rect 1756 215 1896 249
rect 1930 215 1946 249
rect 1576 138 1601 171
rect 1526 105 1601 138
rect 1756 159 1946 215
rect 1756 125 1896 159
rect 1930 125 1946 159
rect 1756 113 1946 125
rect 1277 53 1490 87
rect 1756 79 1762 113
rect 1796 79 1834 113
rect 1868 79 1906 113
rect 1940 79 1946 113
rect 2036 221 2052 255
rect 2086 221 2102 255
rect 2036 155 2102 221
rect 2036 121 2052 155
rect 2086 121 2102 155
rect 2036 105 2102 121
rect 2138 283 2256 299
rect 2138 249 2172 283
rect 2206 249 2256 283
rect 2138 183 2256 249
rect 2138 149 2172 183
rect 2206 149 2256 183
rect 2138 113 2256 149
rect 2328 279 2378 437
rect 2362 245 2378 279
rect 2328 187 2378 245
rect 2362 153 2378 187
rect 2328 137 2378 153
rect 1756 73 1946 79
rect 2138 79 2144 113
rect 2178 79 2216 113
rect 2250 79 2256 113
rect 2138 73 2256 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 114 701 148 735
rect 186 701 220 735
rect 258 701 292 735
rect 450 701 484 735
rect 1020 703 1054 737
rect 1092 703 1126 737
rect 1164 731 1198 737
rect 1164 703 1188 731
rect 1188 703 1198 731
rect 118 79 152 113
rect 190 79 224 113
rect 262 79 296 113
rect 443 79 477 113
rect 515 79 549 113
rect 1769 701 1803 735
rect 1841 701 1875 735
rect 1913 731 1947 735
rect 1913 701 1937 731
rect 1937 701 1947 731
rect 1057 79 1091 113
rect 1129 79 1163 113
rect 1201 79 1235 113
rect 2151 731 2185 735
rect 2151 701 2172 731
rect 2172 701 2185 731
rect 2223 701 2257 735
rect 1762 79 1796 113
rect 1834 79 1868 113
rect 1906 79 1940 113
rect 2144 79 2178 113
rect 2216 79 2250 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 831 2400 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2400 831
rect 0 791 2400 797
rect 0 737 2400 763
rect 0 735 1020 737
rect 0 701 114 735
rect 148 701 186 735
rect 220 701 258 735
rect 292 701 450 735
rect 484 703 1020 735
rect 1054 703 1092 737
rect 1126 703 1164 737
rect 1198 735 2400 737
rect 1198 703 1769 735
rect 484 701 1769 703
rect 1803 701 1841 735
rect 1875 701 1913 735
rect 1947 701 2151 735
rect 2185 701 2223 735
rect 2257 701 2400 735
rect 0 689 2400 701
rect 0 113 2400 125
rect 0 79 118 113
rect 152 79 190 113
rect 224 79 262 113
rect 296 79 443 113
rect 477 79 515 113
rect 549 79 1057 113
rect 1091 79 1129 113
rect 1163 79 1201 113
rect 1235 79 1762 113
rect 1796 79 1834 113
rect 1868 79 1906 113
rect 1940 79 2144 113
rect 2178 79 2216 113
rect 2250 79 2400 113
rect 0 51 2400 79
rect 0 17 2400 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -23 2400 -17
<< labels >>
flabel comment s 831 373 831 373 0 FreeSans 200 90 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfxtp_1
flabel metal1 s 0 51 2400 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 2400 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 689 2400 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 791 2400 814 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2335 168 2369 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2335 242 2369 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2335 316 2369 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2335 390 2369 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2335 464 2369 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2335 538 2369 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2335 612 2369 646 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2400 814
string GDS_END 1154778
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1130742
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
