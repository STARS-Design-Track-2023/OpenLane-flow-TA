magic
tech sky130A
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_0
timestamp 1686671242
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_1
timestamp 1686671242
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_0
timestamp 1686671242
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_1
timestamp 1686671242
transform 1 0 412 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 8131894
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8129944
<< end >>
