magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 98 157 638 203
rect 1 21 638 157
rect 30 -17 64 21
<< locali >>
rect 17 199 66 323
rect 470 119 536 425
rect 570 153 627 323
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 391 69 493
rect 103 425 175 527
rect 17 357 175 391
rect 100 265 175 357
rect 209 345 257 493
rect 291 379 357 527
rect 397 459 627 493
rect 397 345 431 459
rect 209 311 431 345
rect 100 199 436 265
rect 100 165 175 199
rect 17 131 175 165
rect 209 131 436 165
rect 17 51 69 131
rect 103 17 175 97
rect 209 51 248 131
rect 282 17 354 97
rect 388 85 436 131
rect 570 357 627 459
rect 570 85 627 119
rect 388 51 627 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 570 153 627 323 6 A
port 1 nsew signal input
rlabel locali s 17 199 66 323 6 TE
port 2 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 638 157 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 98 157 638 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 470 119 536 425 6 Z
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2030880
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2024692
<< end >>
