magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 992 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 267 47 297 177
rect 351 47 381 177
rect 435 47 465 177
rect 519 47 549 177
rect 606 47 636 177
rect 690 47 720 177
rect 774 47 804 177
rect 858 47 888 177
<< scpmoshvt >>
rect 79 297 109 497
rect 267 297 297 497
rect 351 297 381 497
rect 435 297 465 497
rect 519 297 549 497
rect 606 297 636 497
rect 690 297 720 497
rect 774 297 804 497
rect 858 297 888 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 93 161 177
rect 109 59 119 93
rect 153 59 161 93
rect 109 47 161 59
rect 215 161 267 177
rect 215 127 223 161
rect 257 127 267 161
rect 215 93 267 127
rect 215 59 223 93
rect 257 59 267 93
rect 215 47 267 59
rect 297 161 351 177
rect 297 127 307 161
rect 341 127 351 161
rect 297 47 351 127
rect 381 93 435 177
rect 381 59 391 93
rect 425 59 435 93
rect 381 47 435 59
rect 465 161 519 177
rect 465 127 475 161
rect 509 127 519 161
rect 465 47 519 127
rect 549 161 606 177
rect 549 127 562 161
rect 596 127 606 161
rect 549 93 606 127
rect 549 59 562 93
rect 596 59 606 93
rect 549 47 606 59
rect 636 93 690 177
rect 636 59 646 93
rect 680 59 690 93
rect 636 47 690 59
rect 720 161 774 177
rect 720 127 730 161
rect 764 127 774 161
rect 720 93 774 127
rect 720 59 730 93
rect 764 59 774 93
rect 720 47 774 59
rect 804 93 858 177
rect 804 59 814 93
rect 848 59 858 93
rect 804 47 858 59
rect 888 161 966 177
rect 888 127 920 161
rect 954 127 966 161
rect 888 93 966 127
rect 888 59 920 93
rect 954 59 966 93
rect 888 47 966 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 161 497
rect 109 451 119 485
rect 153 451 161 485
rect 109 417 161 451
rect 109 383 119 417
rect 153 383 161 417
rect 109 297 161 383
rect 215 485 267 497
rect 215 451 223 485
rect 257 451 267 485
rect 215 417 267 451
rect 215 383 223 417
rect 257 383 267 417
rect 215 349 267 383
rect 215 315 223 349
rect 257 315 267 349
rect 215 297 267 315
rect 297 485 351 497
rect 297 451 307 485
rect 341 451 351 485
rect 297 417 351 451
rect 297 383 307 417
rect 341 383 351 417
rect 297 349 351 383
rect 297 315 307 349
rect 341 315 351 349
rect 297 297 351 315
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 297 435 383
rect 465 485 519 497
rect 465 451 475 485
rect 509 451 519 485
rect 465 417 519 451
rect 465 383 475 417
rect 509 383 519 417
rect 465 349 519 383
rect 465 315 475 349
rect 509 315 519 349
rect 465 297 519 315
rect 549 485 606 497
rect 549 451 562 485
rect 596 451 606 485
rect 549 417 606 451
rect 549 383 562 417
rect 596 383 606 417
rect 549 297 606 383
rect 636 485 690 497
rect 636 451 646 485
rect 680 451 690 485
rect 636 417 690 451
rect 636 383 646 417
rect 680 383 690 417
rect 636 349 690 383
rect 636 315 646 349
rect 680 315 690 349
rect 636 297 690 315
rect 720 485 774 497
rect 720 451 730 485
rect 764 451 774 485
rect 720 417 774 451
rect 720 383 730 417
rect 764 383 774 417
rect 720 297 774 383
rect 804 485 858 497
rect 804 451 814 485
rect 848 451 858 485
rect 804 417 858 451
rect 804 383 814 417
rect 848 383 858 417
rect 804 349 858 383
rect 804 315 814 349
rect 848 315 858 349
rect 804 297 858 315
rect 888 485 966 497
rect 888 451 920 485
rect 954 451 966 485
rect 888 417 966 451
rect 888 383 920 417
rect 954 383 966 417
rect 888 349 966 383
rect 888 315 920 349
rect 954 315 966 349
rect 888 297 966 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 59 153 93
rect 223 127 257 161
rect 223 59 257 93
rect 307 127 341 161
rect 391 59 425 93
rect 475 127 509 161
rect 562 127 596 161
rect 562 59 596 93
rect 646 59 680 93
rect 730 127 764 161
rect 730 59 764 93
rect 814 59 848 93
rect 920 127 954 161
rect 920 59 954 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 223 451 257 485
rect 223 383 257 417
rect 223 315 257 349
rect 307 451 341 485
rect 307 383 341 417
rect 307 315 341 349
rect 391 451 425 485
rect 391 383 425 417
rect 475 451 509 485
rect 475 383 509 417
rect 475 315 509 349
rect 562 451 596 485
rect 562 383 596 417
rect 646 451 680 485
rect 646 383 680 417
rect 646 315 680 349
rect 730 451 764 485
rect 730 383 764 417
rect 814 451 848 485
rect 814 383 848 417
rect 814 315 848 349
rect 920 451 954 485
rect 920 383 954 417
rect 920 315 954 349
<< poly >>
rect 79 497 109 523
rect 267 497 297 523
rect 351 497 381 523
rect 435 497 465 523
rect 519 497 549 523
rect 606 497 636 523
rect 690 497 720 523
rect 774 497 804 523
rect 858 497 888 523
rect 79 261 109 297
rect 22 249 109 261
rect 267 259 297 297
rect 351 259 381 297
rect 435 259 465 297
rect 519 259 549 297
rect 22 215 38 249
rect 72 215 109 249
rect 22 203 109 215
rect 201 249 549 259
rect 201 215 217 249
rect 251 215 307 249
rect 341 215 391 249
rect 425 215 549 249
rect 201 205 549 215
rect 79 177 109 203
rect 267 177 297 205
rect 351 177 381 205
rect 435 177 465 205
rect 519 177 549 205
rect 606 259 636 297
rect 690 259 720 297
rect 774 259 804 297
rect 858 259 888 297
rect 606 249 954 259
rect 606 215 647 249
rect 681 215 730 249
rect 764 215 813 249
rect 847 215 904 249
rect 938 215 954 249
rect 606 205 954 215
rect 606 177 636 205
rect 690 177 720 205
rect 774 177 804 205
rect 858 177 888 205
rect 79 21 109 47
rect 267 21 297 47
rect 351 21 381 47
rect 435 21 465 47
rect 519 21 549 47
rect 606 21 636 47
rect 690 21 720 47
rect 774 21 804 47
rect 858 21 888 47
<< polycont >>
rect 38 215 72 249
rect 217 215 251 249
rect 307 215 341 249
rect 391 215 425 249
rect 647 215 681 249
rect 730 215 764 249
rect 813 215 847 249
rect 904 215 938 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 18 485 85 493
rect 18 451 35 485
rect 69 451 85 485
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 18 349 85 383
rect 119 485 257 527
rect 153 451 223 485
rect 119 417 257 451
rect 153 383 223 417
rect 119 367 257 383
rect 18 315 35 349
rect 69 333 85 349
rect 194 349 257 367
rect 69 315 156 333
rect 18 289 156 315
rect 194 315 223 349
rect 194 289 257 315
rect 291 485 357 493
rect 291 451 307 485
rect 341 451 357 485
rect 291 417 357 451
rect 291 383 307 417
rect 341 383 357 417
rect 291 349 357 383
rect 391 485 425 527
rect 391 417 425 451
rect 391 367 425 383
rect 459 485 528 493
rect 459 451 475 485
rect 509 451 528 485
rect 459 417 528 451
rect 459 383 475 417
rect 509 383 528 417
rect 291 315 307 349
rect 341 333 357 349
rect 459 349 528 383
rect 562 485 596 527
rect 562 417 596 451
rect 562 367 596 383
rect 630 485 696 493
rect 630 451 646 485
rect 680 451 696 485
rect 630 417 696 451
rect 630 383 646 417
rect 680 383 696 417
rect 459 333 475 349
rect 341 315 475 333
rect 509 333 528 349
rect 630 349 696 383
rect 730 485 764 527
rect 730 417 764 451
rect 730 367 764 383
rect 798 485 864 493
rect 798 451 814 485
rect 848 451 864 485
rect 798 417 864 451
rect 798 383 814 417
rect 848 383 864 417
rect 630 333 646 349
rect 509 315 646 333
rect 680 333 696 349
rect 798 349 864 383
rect 798 333 814 349
rect 680 315 814 333
rect 848 315 864 349
rect 291 289 864 315
rect 904 485 970 527
rect 904 451 920 485
rect 954 451 970 485
rect 904 417 970 451
rect 904 383 920 417
rect 954 383 970 417
rect 904 349 970 383
rect 904 315 920 349
rect 954 315 970 349
rect 904 299 970 315
rect 122 255 156 289
rect 22 249 88 255
rect 22 215 38 249
rect 72 215 88 249
rect 122 249 441 255
rect 122 215 217 249
rect 251 215 307 249
rect 341 215 391 249
rect 425 215 441 249
rect 122 181 156 215
rect 475 181 528 289
rect 631 249 988 255
rect 631 215 647 249
rect 681 215 730 249
rect 764 215 813 249
rect 847 215 904 249
rect 938 215 988 249
rect 18 161 156 181
rect 18 127 35 161
rect 69 143 156 161
rect 207 161 257 181
rect 69 127 85 143
rect 18 93 85 127
rect 207 127 223 161
rect 291 161 528 181
rect 291 127 307 161
rect 341 127 475 161
rect 509 127 528 161
rect 562 161 970 181
rect 596 143 730 161
rect 596 127 612 143
rect 18 59 35 93
rect 69 59 85 93
rect 18 51 85 59
rect 119 93 158 109
rect 153 59 158 93
rect 119 17 158 59
rect 207 93 257 127
rect 562 93 612 127
rect 714 127 730 143
rect 764 143 920 161
rect 764 127 780 143
rect 207 59 223 93
rect 257 59 391 93
rect 425 59 562 93
rect 596 59 612 93
rect 207 51 612 59
rect 646 93 680 109
rect 646 17 680 59
rect 714 93 780 127
rect 904 127 920 143
rect 954 127 970 161
rect 714 59 730 93
rect 764 59 780 93
rect 714 51 780 59
rect 814 93 862 109
rect 848 59 862 93
rect 814 17 862 59
rect 904 93 970 127
rect 904 59 920 93
rect 954 59 970 93
rect 904 51 970 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel locali s 954 221 988 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 862 221 896 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 770 221 804 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 678 221 712 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel locali s 494 153 528 187 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 494 221 528 255 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 494 289 528 323 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand2b_4
rlabel metal1 s 0 -48 1012 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_END 1820282
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1811226
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 25.300 0.000 
<< end >>
