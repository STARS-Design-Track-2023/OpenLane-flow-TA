magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< metal3 >>
rect 2908 38478 4894 38507
rect 2908 34894 2949 38478
rect 4853 34894 4894 38478
rect 2908 34866 4894 34894
rect 5280 38483 7266 38507
rect 5280 34899 5321 38483
rect 7225 34899 7266 38483
rect 5280 34876 7266 34899
rect 7624 18529 9746 18550
rect 7624 13665 7653 18529
rect 9717 13665 9746 18529
rect 7624 13644 9746 13665
rect 5216 5618 7336 5660
rect 5216 4834 5244 5618
rect 7308 4834 7336 5618
rect 5216 4792 7336 4834
rect 7604 4409 9750 4450
rect 7604 3625 7645 4409
rect 9709 3625 9750 4409
rect 7604 3584 9750 3625
<< via3 >>
rect 2949 34894 4853 38478
rect 5321 34899 7225 38483
rect 7653 13665 9717 18529
rect 5244 4834 7308 5618
rect 7645 3625 9709 4409
<< metal4 >>
rect 2908 38478 4894 38501
rect 2908 34894 2949 38478
rect 4853 34894 4894 38478
rect 2908 34866 4894 34894
rect 5280 38483 7266 38501
rect 5280 34899 5321 38483
rect 7225 34899 7266 38483
rect 5280 34876 7266 34899
rect 7624 18529 9746 18550
rect 7624 13665 7653 18529
rect 9717 13665 9746 18529
rect 7624 13644 9746 13665
rect 5216 5618 7336 5660
rect 5216 4834 5244 5618
rect 7308 4834 7336 5618
rect 5216 4792 7336 4834
rect 7604 4409 9750 4450
rect 7604 3625 7645 4409
rect 9709 3625 9750 4409
rect 7604 3584 9750 3625
<< properties >>
string FIXED_BBOX 0 -406 15000 39592
string GDS_END 2675870
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 2402138
<< end >>
