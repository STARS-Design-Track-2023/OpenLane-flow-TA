magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< pwell >>
rect 894 821 918 872
<< obsli1 >>
rect 0 0 1716 1568
<< obsm1 >>
rect 0 1502 1716 1568
rect 0 66 66 1502
rect 99 816 127 1474
rect 155 844 183 1502
rect 211 816 239 1474
rect 267 844 295 1502
rect 323 816 351 1474
rect 379 844 407 1502
rect 435 816 463 1474
rect 491 844 519 1502
rect 547 816 575 1474
rect 603 844 631 1502
rect 659 816 687 1474
rect 715 844 743 1502
rect 771 816 799 1474
rect 831 816 885 1474
rect 917 816 945 1474
rect 973 844 1001 1502
rect 1029 816 1057 1474
rect 1085 844 1113 1502
rect 1141 816 1169 1474
rect 1197 844 1225 1502
rect 1253 816 1281 1474
rect 1309 844 1337 1502
rect 1365 816 1393 1474
rect 1421 844 1449 1502
rect 1477 816 1505 1474
rect 1533 844 1561 1502
rect 1589 816 1617 1474
rect 99 752 1617 816
rect 99 94 127 752
rect 155 66 183 724
rect 211 94 239 752
rect 267 66 295 724
rect 323 94 351 752
rect 379 66 407 724
rect 435 94 463 752
rect 491 66 519 724
rect 547 94 575 752
rect 603 66 631 724
rect 659 94 687 752
rect 715 66 743 724
rect 771 94 799 752
rect 831 94 885 752
rect 917 94 945 752
rect 973 66 1001 724
rect 1029 94 1057 752
rect 1085 66 1113 724
rect 1141 94 1169 752
rect 1197 66 1225 724
rect 1253 94 1281 752
rect 1309 66 1337 724
rect 1365 94 1393 752
rect 1421 66 1449 724
rect 1477 94 1505 752
rect 1533 66 1561 724
rect 1589 94 1617 752
rect 1650 66 1716 1502
rect 0 0 1716 66
<< obsm2 >>
rect 0 1502 803 1568
rect 0 1418 66 1502
rect 831 1474 885 1568
rect 913 1502 1716 1568
rect 94 1446 1622 1474
rect 0 1390 802 1418
rect 0 1306 66 1390
rect 830 1362 886 1446
rect 1650 1418 1716 1502
rect 914 1390 1716 1418
rect 94 1334 1622 1362
rect 0 1278 802 1306
rect 0 1194 66 1278
rect 830 1250 886 1334
rect 1650 1306 1716 1390
rect 914 1278 1716 1306
rect 94 1222 1622 1250
rect 0 1166 802 1194
rect 0 1082 66 1166
rect 830 1138 886 1222
rect 1650 1194 1716 1278
rect 914 1166 1716 1194
rect 94 1110 1622 1138
rect 0 1054 802 1082
rect 0 970 66 1054
rect 830 1026 886 1110
rect 1650 1082 1716 1166
rect 914 1054 1716 1082
rect 94 998 1622 1026
rect 0 942 802 970
rect 0 839 66 942
rect 830 914 886 998
rect 1650 970 1716 1054
rect 914 942 1716 970
rect 94 840 1622 914
rect 830 812 886 840
rect 1650 839 1716 942
rect 74 811 1642 812
rect 0 757 1716 811
rect 74 756 1642 757
rect 0 626 66 729
rect 830 728 886 756
rect 94 654 1622 728
rect 0 598 802 626
rect 0 514 66 598
rect 830 570 886 654
rect 1650 626 1716 729
rect 914 598 1716 626
rect 94 542 1622 570
rect 0 486 802 514
rect 0 402 66 486
rect 830 458 886 542
rect 1650 514 1716 598
rect 914 486 1716 514
rect 94 430 1622 458
rect 0 374 802 402
rect 0 290 66 374
rect 830 346 886 430
rect 1650 402 1716 486
rect 914 374 1716 402
rect 94 318 1622 346
rect 0 262 802 290
rect 0 178 66 262
rect 830 234 886 318
rect 1650 290 1716 374
rect 914 262 1716 290
rect 94 206 1622 234
rect 0 150 802 178
rect 0 66 66 150
rect 830 122 886 206
rect 1650 178 1716 262
rect 914 150 1716 178
rect 94 94 1622 122
rect 0 0 803 66
rect 831 0 885 94
rect 1650 66 1716 150
rect 913 0 1716 66
<< metal3 >>
rect 0 1502 1716 1568
rect 0 66 66 1502
rect 126 817 204 1442
rect 264 877 342 1502
rect 402 817 480 1442
rect 540 877 618 1502
rect 678 817 756 1442
rect 819 877 897 1502
rect 960 817 1038 1442
rect 1098 877 1176 1502
rect 1236 817 1314 1442
rect 1374 877 1452 1502
rect 1512 817 1590 1442
rect 126 751 1590 817
rect 126 126 204 751
rect 264 66 342 691
rect 402 126 480 751
rect 540 66 618 691
rect 678 126 756 751
rect 819 66 897 691
rect 960 126 1038 751
rect 1098 66 1176 691
rect 1236 126 1314 751
rect 1374 66 1452 691
rect 1512 126 1590 751
rect 1650 66 1716 1502
rect 0 0 1716 66
<< obsm4 >>
rect 63 1103 465 1505
rect 658 1103 1060 1505
rect 1251 1103 1653 1505
rect 63 584 465 986
rect 658 584 1060 986
rect 1251 584 1653 986
rect 63 63 465 465
rect 658 63 1060 465
rect 1251 63 1653 465
<< metal5 >>
rect 0 0 1716 1568
<< labels >>
rlabel metal3 s 1650 66 1716 1502 6 C0
port 1 nsew
rlabel metal3 s 1374 877 1452 1502 6 C0
port 1 nsew
rlabel metal3 s 1374 66 1452 691 6 C0
port 1 nsew
rlabel metal3 s 1098 877 1176 1502 6 C0
port 1 nsew
rlabel metal3 s 1098 66 1176 691 6 C0
port 1 nsew
rlabel metal3 s 819 877 897 1502 6 C0
port 1 nsew
rlabel metal3 s 819 66 897 691 6 C0
port 1 nsew
rlabel metal3 s 540 877 618 1502 6 C0
port 1 nsew
rlabel metal3 s 540 66 618 691 6 C0
port 1 nsew
rlabel metal3 s 264 877 342 1502 6 C0
port 1 nsew
rlabel metal3 s 264 66 342 691 6 C0
port 1 nsew
rlabel metal3 s 0 1502 1716 1568 6 C0
port 1 nsew
rlabel metal3 s 0 66 66 1502 6 C0
port 1 nsew
rlabel metal3 s 0 0 1716 66 6 C0
port 1 nsew
rlabel metal3 s 1512 817 1590 1442 6 C1
port 2 nsew
rlabel metal3 s 1512 126 1590 751 6 C1
port 2 nsew
rlabel metal3 s 1236 817 1314 1442 6 C1
port 2 nsew
rlabel metal3 s 1236 126 1314 751 6 C1
port 2 nsew
rlabel metal3 s 960 817 1038 1442 6 C1
port 2 nsew
rlabel metal3 s 960 126 1038 751 6 C1
port 2 nsew
rlabel metal3 s 678 817 756 1442 6 C1
port 2 nsew
rlabel metal3 s 678 126 756 751 6 C1
port 2 nsew
rlabel metal3 s 402 817 480 1442 6 C1
port 2 nsew
rlabel metal3 s 402 126 480 751 6 C1
port 2 nsew
rlabel metal3 s 126 817 204 1442 6 C1
port 2 nsew
rlabel metal3 s 126 751 1590 817 6 C1
port 2 nsew
rlabel metal3 s 126 126 204 751 6 C1
port 2 nsew
rlabel metal5 s 0 0 1716 1568 6 MET5
port 4 nsew
rlabel pwell s 894 821 918 872 6 SUB
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1716 1568
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 534570
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 506342
string device primitive
<< end >>
