magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__hvdfm1sd2__example_55959141808719  sky130_fd_pr__hvdfm1sd2__example_55959141808719_0
timestamp 1686671242
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808782  sky130_fd_pr__hvdfm1sd__example_55959141808782_0
timestamp 1686671242
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 27736648
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 27735592
<< end >>
