magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_0
timestamp 1686671242
transform -1 0 -7 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_1
timestamp 1686671242
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_2
timestamp 1686671242
transform 1 0 263 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_3
timestamp 1686671242
transform 1 0 426 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_4
timestamp 1686671242
transform 1 0 589 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_5
timestamp 1686671242
transform 1 0 752 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_6
timestamp 1686671242
transform 1 0 915 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 8673962
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8669930
<< end >>
