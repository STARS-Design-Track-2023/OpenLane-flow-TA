magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< pwell >>
rect 1176 1289 1197 1338
<< metal1 >>
rect 0 2331 2282 2338
rect 0 2282 88 2331
rect 0 2230 7 2282
rect 59 2279 88 2282
rect 140 2279 152 2331
rect 204 2279 216 2331
rect 268 2279 280 2331
rect 332 2279 344 2331
rect 396 2279 408 2331
rect 460 2279 472 2331
rect 524 2279 536 2331
rect 588 2279 600 2331
rect 652 2279 664 2331
rect 716 2279 728 2331
rect 780 2279 792 2331
rect 844 2279 856 2331
rect 908 2279 920 2331
rect 972 2279 984 2331
rect 1036 2279 1246 2331
rect 1298 2279 1310 2331
rect 1362 2279 1374 2331
rect 1426 2279 1438 2331
rect 1490 2279 1502 2331
rect 1554 2279 1566 2331
rect 1618 2279 1630 2331
rect 1682 2279 1694 2331
rect 1746 2279 1758 2331
rect 1810 2279 1822 2331
rect 1874 2279 1886 2331
rect 1938 2279 1950 2331
rect 2002 2279 2014 2331
rect 2066 2279 2078 2331
rect 2130 2279 2142 2331
rect 2194 2282 2282 2331
rect 2194 2279 2223 2282
rect 59 2272 2223 2279
rect 59 2230 72 2272
rect 0 2218 72 2230
rect 0 2166 7 2218
rect 59 2166 72 2218
rect 0 2154 72 2166
rect 0 2102 7 2154
rect 59 2102 72 2154
rect 0 2090 72 2102
rect 0 2038 7 2090
rect 59 2038 72 2090
rect 0 2026 72 2038
rect 0 1974 7 2026
rect 59 1974 72 2026
rect 0 1962 72 1974
rect 0 1910 7 1962
rect 59 1910 72 1962
rect 0 1898 72 1910
rect 0 1846 7 1898
rect 59 1846 72 1898
rect 0 1834 72 1846
rect 0 1782 7 1834
rect 59 1782 72 1834
rect 0 1770 72 1782
rect 0 1718 7 1770
rect 59 1718 72 1770
rect 0 1706 72 1718
rect 0 1654 7 1706
rect 59 1654 72 1706
rect 0 1642 72 1654
rect 0 1590 7 1642
rect 59 1590 72 1642
rect 0 1578 72 1590
rect 0 1526 7 1578
rect 59 1526 72 1578
rect 0 1514 72 1526
rect 0 1462 7 1514
rect 59 1462 72 1514
rect 0 1450 72 1462
rect 0 1398 7 1450
rect 59 1398 72 1450
rect 0 1386 72 1398
rect 0 1334 7 1386
rect 59 1334 72 1386
rect 0 1322 72 1334
rect 0 1270 7 1322
rect 59 1270 72 1322
rect 0 1068 72 1270
rect 0 1016 7 1068
rect 59 1016 72 1068
rect 0 1004 72 1016
rect 0 952 7 1004
rect 59 952 72 1004
rect 0 940 72 952
rect 0 888 7 940
rect 59 888 72 940
rect 0 876 72 888
rect 0 824 7 876
rect 59 824 72 876
rect 0 812 72 824
rect 0 760 7 812
rect 59 760 72 812
rect 0 748 72 760
rect 0 696 7 748
rect 59 696 72 748
rect 0 684 72 696
rect 0 632 7 684
rect 59 632 72 684
rect 0 620 72 632
rect 0 568 7 620
rect 59 568 72 620
rect 0 556 72 568
rect 0 504 7 556
rect 59 504 72 556
rect 0 492 72 504
rect 0 440 7 492
rect 59 440 72 492
rect 0 428 72 440
rect 0 376 7 428
rect 59 376 72 428
rect 0 364 72 376
rect 0 312 7 364
rect 59 312 72 364
rect 0 300 72 312
rect 0 248 7 300
rect 59 248 72 300
rect 0 236 72 248
rect 0 184 7 236
rect 59 184 72 236
rect 0 172 72 184
rect 0 120 7 172
rect 59 120 72 172
rect 0 108 72 120
rect 0 56 7 108
rect 59 66 72 108
rect 100 1201 128 2244
rect 156 1229 184 2272
rect 212 1201 240 2244
rect 268 1229 296 2272
rect 324 1201 352 2244
rect 380 1229 408 2272
rect 436 1201 464 2244
rect 492 1229 520 2272
rect 548 1201 576 2244
rect 604 1229 632 2272
rect 660 1201 688 2244
rect 716 1229 744 2272
rect 772 1201 800 2244
rect 828 1229 856 2272
rect 884 1201 912 2244
rect 940 1229 968 2272
rect 996 1201 1024 2244
rect 1052 1229 1080 2272
rect 1108 2237 1174 2244
rect 1108 2185 1115 2237
rect 1167 2185 1174 2237
rect 1108 2173 1174 2185
rect 1108 2121 1115 2173
rect 1167 2121 1174 2173
rect 1108 2109 1174 2121
rect 1108 2057 1115 2109
rect 1167 2057 1174 2109
rect 1108 2045 1174 2057
rect 1108 1993 1115 2045
rect 1167 1993 1174 2045
rect 1108 1981 1174 1993
rect 1108 1929 1115 1981
rect 1167 1929 1174 1981
rect 1108 1917 1174 1929
rect 1108 1865 1115 1917
rect 1167 1865 1174 1917
rect 1108 1853 1174 1865
rect 1108 1801 1115 1853
rect 1167 1801 1174 1853
rect 1108 1789 1174 1801
rect 1108 1737 1115 1789
rect 1167 1737 1174 1789
rect 1108 1725 1174 1737
rect 1108 1673 1115 1725
rect 1167 1673 1174 1725
rect 1108 1661 1174 1673
rect 1108 1609 1115 1661
rect 1167 1609 1174 1661
rect 1108 1597 1174 1609
rect 1108 1545 1115 1597
rect 1167 1545 1174 1597
rect 1108 1533 1174 1545
rect 1108 1481 1115 1533
rect 1167 1481 1174 1533
rect 1108 1469 1174 1481
rect 1108 1417 1115 1469
rect 1167 1417 1174 1469
rect 1108 1405 1174 1417
rect 1108 1353 1115 1405
rect 1167 1353 1174 1405
rect 1108 1341 1174 1353
rect 1108 1289 1115 1341
rect 1167 1289 1174 1341
rect 1108 1277 1174 1289
rect 1108 1225 1115 1277
rect 1167 1225 1174 1277
rect 1202 1229 1230 2272
rect 1108 1201 1174 1225
rect 1258 1201 1286 2244
rect 1314 1229 1342 2272
rect 1370 1201 1398 2244
rect 1426 1229 1454 2272
rect 1482 1201 1510 2244
rect 1538 1229 1566 2272
rect 1594 1201 1622 2244
rect 1650 1229 1678 2272
rect 1706 1201 1734 2244
rect 1762 1229 1790 2272
rect 1818 1201 1846 2244
rect 1874 1229 1902 2272
rect 1930 1201 1958 2244
rect 1986 1229 2014 2272
rect 2042 1201 2070 2244
rect 2098 1229 2126 2272
rect 2154 1201 2182 2244
rect 100 1195 2182 1201
rect 100 1143 152 1195
rect 204 1143 216 1195
rect 268 1143 280 1195
rect 332 1143 344 1195
rect 396 1143 408 1195
rect 460 1143 472 1195
rect 524 1143 536 1195
rect 588 1143 600 1195
rect 652 1143 664 1195
rect 716 1143 728 1195
rect 780 1143 792 1195
rect 844 1143 856 1195
rect 908 1143 920 1195
rect 972 1143 984 1195
rect 1036 1143 1048 1195
rect 1100 1143 1182 1195
rect 1234 1143 1246 1195
rect 1298 1143 1310 1195
rect 1362 1143 1374 1195
rect 1426 1143 1438 1195
rect 1490 1143 1502 1195
rect 1554 1143 1566 1195
rect 1618 1143 1630 1195
rect 1682 1143 1694 1195
rect 1746 1143 1758 1195
rect 1810 1143 1822 1195
rect 1874 1143 1886 1195
rect 1938 1143 1950 1195
rect 2002 1143 2014 1195
rect 2066 1143 2078 1195
rect 2130 1143 2182 1195
rect 100 1137 2182 1143
rect 100 94 128 1137
rect 156 66 184 1109
rect 212 94 240 1137
rect 268 66 296 1109
rect 324 94 352 1137
rect 380 66 408 1109
rect 436 94 464 1137
rect 492 66 520 1109
rect 548 94 576 1137
rect 604 66 632 1109
rect 660 94 688 1137
rect 716 66 744 1109
rect 772 94 800 1137
rect 828 66 856 1109
rect 884 94 912 1137
rect 940 66 968 1109
rect 996 94 1024 1137
rect 1108 1113 1174 1137
rect 1052 66 1080 1109
rect 1108 1061 1115 1113
rect 1167 1061 1174 1113
rect 1108 1049 1174 1061
rect 1108 997 1115 1049
rect 1167 997 1174 1049
rect 1108 985 1174 997
rect 1108 933 1115 985
rect 1167 933 1174 985
rect 1108 921 1174 933
rect 1108 869 1115 921
rect 1167 869 1174 921
rect 1108 857 1174 869
rect 1108 805 1115 857
rect 1167 805 1174 857
rect 1108 793 1174 805
rect 1108 741 1115 793
rect 1167 741 1174 793
rect 1108 729 1174 741
rect 1108 677 1115 729
rect 1167 677 1174 729
rect 1108 665 1174 677
rect 1108 613 1115 665
rect 1167 613 1174 665
rect 1108 601 1174 613
rect 1108 549 1115 601
rect 1167 549 1174 601
rect 1108 537 1174 549
rect 1108 485 1115 537
rect 1167 485 1174 537
rect 1108 473 1174 485
rect 1108 421 1115 473
rect 1167 421 1174 473
rect 1108 409 1174 421
rect 1108 357 1115 409
rect 1167 357 1174 409
rect 1108 345 1174 357
rect 1108 293 1115 345
rect 1167 293 1174 345
rect 1108 281 1174 293
rect 1108 229 1115 281
rect 1167 229 1174 281
rect 1108 217 1174 229
rect 1108 165 1115 217
rect 1167 165 1174 217
rect 1108 153 1174 165
rect 1108 101 1115 153
rect 1167 101 1174 153
rect 1108 94 1174 101
rect 1202 66 1230 1109
rect 1258 94 1286 1137
rect 1314 66 1342 1109
rect 1370 94 1398 1137
rect 1426 66 1454 1109
rect 1482 94 1510 1137
rect 1538 66 1566 1109
rect 1594 94 1622 1137
rect 1650 66 1678 1109
rect 1706 94 1734 1137
rect 1762 66 1790 1109
rect 1818 94 1846 1137
rect 1874 66 1902 1109
rect 1930 94 1958 1137
rect 1986 66 2014 1109
rect 2042 94 2070 1137
rect 2098 66 2126 1109
rect 2154 94 2182 1137
rect 2210 2230 2223 2272
rect 2275 2230 2282 2282
rect 2210 2218 2282 2230
rect 2210 2166 2223 2218
rect 2275 2166 2282 2218
rect 2210 2154 2282 2166
rect 2210 2102 2223 2154
rect 2275 2102 2282 2154
rect 2210 2090 2282 2102
rect 2210 2038 2223 2090
rect 2275 2038 2282 2090
rect 2210 2026 2282 2038
rect 2210 1974 2223 2026
rect 2275 1974 2282 2026
rect 2210 1962 2282 1974
rect 2210 1910 2223 1962
rect 2275 1910 2282 1962
rect 2210 1898 2282 1910
rect 2210 1846 2223 1898
rect 2275 1846 2282 1898
rect 2210 1834 2282 1846
rect 2210 1782 2223 1834
rect 2275 1782 2282 1834
rect 2210 1770 2282 1782
rect 2210 1718 2223 1770
rect 2275 1718 2282 1770
rect 2210 1706 2282 1718
rect 2210 1654 2223 1706
rect 2275 1654 2282 1706
rect 2210 1642 2282 1654
rect 2210 1590 2223 1642
rect 2275 1590 2282 1642
rect 2210 1578 2282 1590
rect 2210 1526 2223 1578
rect 2275 1526 2282 1578
rect 2210 1514 2282 1526
rect 2210 1462 2223 1514
rect 2275 1462 2282 1514
rect 2210 1450 2282 1462
rect 2210 1398 2223 1450
rect 2275 1398 2282 1450
rect 2210 1386 2282 1398
rect 2210 1334 2223 1386
rect 2275 1334 2282 1386
rect 2210 1322 2282 1334
rect 2210 1270 2223 1322
rect 2275 1270 2282 1322
rect 2210 1068 2282 1270
rect 2210 1016 2223 1068
rect 2275 1016 2282 1068
rect 2210 1004 2282 1016
rect 2210 952 2223 1004
rect 2275 952 2282 1004
rect 2210 940 2282 952
rect 2210 888 2223 940
rect 2275 888 2282 940
rect 2210 876 2282 888
rect 2210 824 2223 876
rect 2275 824 2282 876
rect 2210 812 2282 824
rect 2210 760 2223 812
rect 2275 760 2282 812
rect 2210 748 2282 760
rect 2210 696 2223 748
rect 2275 696 2282 748
rect 2210 684 2282 696
rect 2210 632 2223 684
rect 2275 632 2282 684
rect 2210 620 2282 632
rect 2210 568 2223 620
rect 2275 568 2282 620
rect 2210 556 2282 568
rect 2210 504 2223 556
rect 2275 504 2282 556
rect 2210 492 2282 504
rect 2210 440 2223 492
rect 2275 440 2282 492
rect 2210 428 2282 440
rect 2210 376 2223 428
rect 2275 376 2282 428
rect 2210 364 2282 376
rect 2210 312 2223 364
rect 2275 312 2282 364
rect 2210 300 2282 312
rect 2210 248 2223 300
rect 2275 248 2282 300
rect 2210 236 2282 248
rect 2210 184 2223 236
rect 2275 184 2282 236
rect 2210 172 2282 184
rect 2210 120 2223 172
rect 2275 120 2282 172
rect 2210 108 2282 120
rect 2210 66 2223 108
rect 59 59 2223 66
rect 59 56 88 59
rect 0 7 88 56
rect 140 7 152 59
rect 204 7 216 59
rect 268 7 280 59
rect 332 7 344 59
rect 396 7 408 59
rect 460 7 472 59
rect 524 7 536 59
rect 588 7 600 59
rect 652 7 664 59
rect 716 7 728 59
rect 780 7 792 59
rect 844 7 856 59
rect 908 7 920 59
rect 972 7 984 59
rect 1036 7 1246 59
rect 1298 7 1310 59
rect 1362 7 1374 59
rect 1426 7 1438 59
rect 1490 7 1502 59
rect 1554 7 1566 59
rect 1618 7 1630 59
rect 1682 7 1694 59
rect 1746 7 1758 59
rect 1810 7 1822 59
rect 1874 7 1886 59
rect 1938 7 1950 59
rect 2002 7 2014 59
rect 2066 7 2078 59
rect 2130 7 2142 59
rect 2194 56 2223 59
rect 2275 56 2282 108
rect 2194 7 2282 56
rect 0 0 2282 7
<< via1 >>
rect 7 2230 59 2282
rect 88 2279 140 2331
rect 152 2279 204 2331
rect 216 2279 268 2331
rect 280 2279 332 2331
rect 344 2279 396 2331
rect 408 2279 460 2331
rect 472 2279 524 2331
rect 536 2279 588 2331
rect 600 2279 652 2331
rect 664 2279 716 2331
rect 728 2279 780 2331
rect 792 2279 844 2331
rect 856 2279 908 2331
rect 920 2279 972 2331
rect 984 2279 1036 2331
rect 1246 2279 1298 2331
rect 1310 2279 1362 2331
rect 1374 2279 1426 2331
rect 1438 2279 1490 2331
rect 1502 2279 1554 2331
rect 1566 2279 1618 2331
rect 1630 2279 1682 2331
rect 1694 2279 1746 2331
rect 1758 2279 1810 2331
rect 1822 2279 1874 2331
rect 1886 2279 1938 2331
rect 1950 2279 2002 2331
rect 2014 2279 2066 2331
rect 2078 2279 2130 2331
rect 2142 2279 2194 2331
rect 7 2166 59 2218
rect 7 2102 59 2154
rect 7 2038 59 2090
rect 7 1974 59 2026
rect 7 1910 59 1962
rect 7 1846 59 1898
rect 7 1782 59 1834
rect 7 1718 59 1770
rect 7 1654 59 1706
rect 7 1590 59 1642
rect 7 1526 59 1578
rect 7 1462 59 1514
rect 7 1398 59 1450
rect 7 1334 59 1386
rect 7 1270 59 1322
rect 7 1016 59 1068
rect 7 952 59 1004
rect 7 888 59 940
rect 7 824 59 876
rect 7 760 59 812
rect 7 696 59 748
rect 7 632 59 684
rect 7 568 59 620
rect 7 504 59 556
rect 7 440 59 492
rect 7 376 59 428
rect 7 312 59 364
rect 7 248 59 300
rect 7 184 59 236
rect 7 120 59 172
rect 7 56 59 108
rect 1115 2185 1167 2237
rect 1115 2121 1167 2173
rect 1115 2057 1167 2109
rect 1115 1993 1167 2045
rect 1115 1929 1167 1981
rect 1115 1865 1167 1917
rect 1115 1801 1167 1853
rect 1115 1737 1167 1789
rect 1115 1673 1167 1725
rect 1115 1609 1167 1661
rect 1115 1545 1167 1597
rect 1115 1481 1167 1533
rect 1115 1417 1167 1469
rect 1115 1353 1167 1405
rect 1115 1289 1167 1341
rect 1115 1225 1167 1277
rect 152 1143 204 1195
rect 216 1143 268 1195
rect 280 1143 332 1195
rect 344 1143 396 1195
rect 408 1143 460 1195
rect 472 1143 524 1195
rect 536 1143 588 1195
rect 600 1143 652 1195
rect 664 1143 716 1195
rect 728 1143 780 1195
rect 792 1143 844 1195
rect 856 1143 908 1195
rect 920 1143 972 1195
rect 984 1143 1036 1195
rect 1048 1143 1100 1195
rect 1182 1143 1234 1195
rect 1246 1143 1298 1195
rect 1310 1143 1362 1195
rect 1374 1143 1426 1195
rect 1438 1143 1490 1195
rect 1502 1143 1554 1195
rect 1566 1143 1618 1195
rect 1630 1143 1682 1195
rect 1694 1143 1746 1195
rect 1758 1143 1810 1195
rect 1822 1143 1874 1195
rect 1886 1143 1938 1195
rect 1950 1143 2002 1195
rect 2014 1143 2066 1195
rect 2078 1143 2130 1195
rect 1115 1061 1167 1113
rect 1115 997 1167 1049
rect 1115 933 1167 985
rect 1115 869 1167 921
rect 1115 805 1167 857
rect 1115 741 1167 793
rect 1115 677 1167 729
rect 1115 613 1167 665
rect 1115 549 1167 601
rect 1115 485 1167 537
rect 1115 421 1167 473
rect 1115 357 1167 409
rect 1115 293 1167 345
rect 1115 229 1167 281
rect 1115 165 1167 217
rect 1115 101 1167 153
rect 2223 2230 2275 2282
rect 2223 2166 2275 2218
rect 2223 2102 2275 2154
rect 2223 2038 2275 2090
rect 2223 1974 2275 2026
rect 2223 1910 2275 1962
rect 2223 1846 2275 1898
rect 2223 1782 2275 1834
rect 2223 1718 2275 1770
rect 2223 1654 2275 1706
rect 2223 1590 2275 1642
rect 2223 1526 2275 1578
rect 2223 1462 2275 1514
rect 2223 1398 2275 1450
rect 2223 1334 2275 1386
rect 2223 1270 2275 1322
rect 2223 1016 2275 1068
rect 2223 952 2275 1004
rect 2223 888 2275 940
rect 2223 824 2275 876
rect 2223 760 2275 812
rect 2223 696 2275 748
rect 2223 632 2275 684
rect 2223 568 2275 620
rect 2223 504 2275 556
rect 2223 440 2275 492
rect 2223 376 2275 428
rect 2223 312 2275 364
rect 2223 248 2275 300
rect 2223 184 2275 236
rect 2223 120 2275 172
rect 88 7 140 59
rect 152 7 204 59
rect 216 7 268 59
rect 280 7 332 59
rect 344 7 396 59
rect 408 7 460 59
rect 472 7 524 59
rect 536 7 588 59
rect 600 7 652 59
rect 664 7 716 59
rect 728 7 780 59
rect 792 7 844 59
rect 856 7 908 59
rect 920 7 972 59
rect 984 7 1036 59
rect 1246 7 1298 59
rect 1310 7 1362 59
rect 1374 7 1426 59
rect 1438 7 1490 59
rect 1502 7 1554 59
rect 1566 7 1618 59
rect 1630 7 1682 59
rect 1694 7 1746 59
rect 1758 7 1810 59
rect 1822 7 1874 59
rect 1886 7 1938 59
rect 1950 7 2002 59
rect 2014 7 2066 59
rect 2078 7 2130 59
rect 2142 7 2194 59
rect 2223 56 2275 108
<< metal2 >>
rect 0 2331 1086 2338
rect 0 2282 88 2331
rect 0 2230 7 2282
rect 59 2279 88 2282
rect 140 2279 152 2331
rect 204 2279 216 2331
rect 268 2279 280 2331
rect 332 2279 344 2331
rect 396 2279 408 2331
rect 460 2279 472 2331
rect 524 2279 536 2331
rect 588 2279 600 2331
rect 652 2279 664 2331
rect 716 2279 728 2331
rect 780 2279 792 2331
rect 844 2279 856 2331
rect 908 2279 920 2331
rect 972 2279 984 2331
rect 1036 2279 1086 2331
rect 59 2272 1086 2279
rect 59 2230 66 2272
rect 1114 2244 1168 2338
rect 1196 2331 2282 2338
rect 1196 2279 1246 2331
rect 1298 2279 1310 2331
rect 1362 2279 1374 2331
rect 1426 2279 1438 2331
rect 1490 2279 1502 2331
rect 1554 2279 1566 2331
rect 1618 2279 1630 2331
rect 1682 2279 1694 2331
rect 1746 2279 1758 2331
rect 1810 2279 1822 2331
rect 1874 2279 1886 2331
rect 1938 2279 1950 2331
rect 2002 2279 2014 2331
rect 2066 2279 2078 2331
rect 2130 2279 2142 2331
rect 2194 2282 2282 2331
rect 2194 2279 2223 2282
rect 1196 2272 2223 2279
rect 0 2218 66 2230
rect 0 2166 7 2218
rect 59 2188 66 2218
rect 94 2237 2188 2244
rect 94 2216 1115 2237
rect 59 2166 1085 2188
rect 0 2160 1085 2166
rect 1113 2185 1115 2216
rect 1167 2216 2188 2237
rect 2216 2230 2223 2272
rect 2275 2230 2282 2282
rect 2216 2218 2282 2230
rect 1167 2185 1169 2216
rect 2216 2188 2223 2218
rect 1113 2173 1169 2185
rect 0 2154 66 2160
rect 0 2102 7 2154
rect 59 2102 66 2154
rect 1113 2132 1115 2173
rect 94 2121 1115 2132
rect 1167 2132 1169 2173
rect 1197 2166 2223 2188
rect 2275 2166 2282 2218
rect 1197 2160 2282 2166
rect 2216 2154 2282 2160
rect 1167 2121 2188 2132
rect 94 2109 2188 2121
rect 94 2104 1115 2109
rect 0 2090 66 2102
rect 0 2038 7 2090
rect 59 2076 66 2090
rect 59 2048 1085 2076
rect 1113 2057 1115 2104
rect 1167 2104 2188 2109
rect 1167 2057 1169 2104
rect 2216 2102 2223 2154
rect 2275 2102 2282 2154
rect 2216 2090 2282 2102
rect 2216 2076 2223 2090
rect 59 2038 66 2048
rect 0 2026 66 2038
rect 0 1974 7 2026
rect 59 1974 66 2026
rect 1113 2045 1169 2057
rect 1197 2048 2223 2076
rect 1113 2020 1115 2045
rect 94 1993 1115 2020
rect 1167 2020 1169 2045
rect 2216 2038 2223 2048
rect 2275 2038 2282 2090
rect 2216 2026 2282 2038
rect 1167 1993 2188 2020
rect 94 1992 2188 1993
rect 0 1964 66 1974
rect 1113 1981 1169 1992
rect 0 1962 1085 1964
rect 0 1910 7 1962
rect 59 1936 1085 1962
rect 59 1910 66 1936
rect 0 1898 66 1910
rect 1113 1929 1115 1981
rect 1167 1929 1169 1981
rect 2216 1974 2223 2026
rect 2275 1974 2282 2026
rect 2216 1964 2282 1974
rect 1197 1962 2282 1964
rect 1197 1936 2223 1962
rect 1113 1917 1169 1929
rect 1113 1908 1115 1917
rect 0 1846 7 1898
rect 59 1852 66 1898
rect 94 1880 1115 1908
rect 1113 1865 1115 1880
rect 1167 1908 1169 1917
rect 2216 1910 2223 1936
rect 2275 1910 2282 1962
rect 1167 1880 2188 1908
rect 2216 1898 2282 1910
rect 1167 1865 1169 1880
rect 1113 1853 1169 1865
rect 59 1846 1085 1852
rect 0 1834 1085 1846
rect 0 1782 7 1834
rect 59 1824 1085 1834
rect 59 1782 66 1824
rect 1113 1801 1115 1853
rect 1167 1801 1169 1853
rect 2216 1852 2223 1898
rect 1197 1846 2223 1852
rect 2275 1846 2282 1898
rect 1197 1834 2282 1846
rect 1197 1824 2223 1834
rect 1113 1796 1169 1801
rect 0 1770 66 1782
rect 0 1718 7 1770
rect 59 1740 66 1770
rect 94 1789 2188 1796
rect 94 1768 1115 1789
rect 59 1718 1085 1740
rect 0 1712 1085 1718
rect 1113 1737 1115 1768
rect 1167 1768 2188 1789
rect 2216 1782 2223 1824
rect 2275 1782 2282 1834
rect 2216 1770 2282 1782
rect 1167 1737 1169 1768
rect 2216 1740 2223 1770
rect 1113 1725 1169 1737
rect 0 1706 66 1712
rect 0 1654 7 1706
rect 59 1654 66 1706
rect 1113 1684 1115 1725
rect 94 1673 1115 1684
rect 1167 1684 1169 1725
rect 1197 1718 2223 1740
rect 2275 1718 2282 1770
rect 1197 1712 2282 1718
rect 2216 1706 2282 1712
rect 1167 1673 2188 1684
rect 94 1661 2188 1673
rect 94 1656 1115 1661
rect 0 1642 66 1654
rect 0 1590 7 1642
rect 59 1628 66 1642
rect 59 1600 1085 1628
rect 1113 1609 1115 1656
rect 1167 1656 2188 1661
rect 1167 1609 1169 1656
rect 2216 1654 2223 1706
rect 2275 1654 2282 1706
rect 2216 1642 2282 1654
rect 2216 1628 2223 1642
rect 59 1590 66 1600
rect 0 1578 66 1590
rect 0 1526 7 1578
rect 59 1526 66 1578
rect 1113 1597 1169 1609
rect 1197 1600 2223 1628
rect 1113 1572 1115 1597
rect 94 1545 1115 1572
rect 1167 1572 1169 1597
rect 2216 1590 2223 1600
rect 2275 1590 2282 1642
rect 2216 1578 2282 1590
rect 1167 1545 2188 1572
rect 94 1544 2188 1545
rect 0 1516 66 1526
rect 1113 1533 1169 1544
rect 0 1514 1085 1516
rect 0 1462 7 1514
rect 59 1488 1085 1514
rect 59 1462 66 1488
rect 0 1450 66 1462
rect 1113 1481 1115 1533
rect 1167 1481 1169 1533
rect 2216 1526 2223 1578
rect 2275 1526 2282 1578
rect 2216 1516 2282 1526
rect 1197 1514 2282 1516
rect 1197 1488 2223 1514
rect 1113 1469 1169 1481
rect 1113 1460 1115 1469
rect 0 1398 7 1450
rect 59 1404 66 1450
rect 94 1432 1115 1460
rect 1113 1417 1115 1432
rect 1167 1460 1169 1469
rect 2216 1462 2223 1488
rect 2275 1462 2282 1514
rect 1167 1432 2188 1460
rect 2216 1450 2282 1462
rect 1167 1417 1169 1432
rect 1113 1405 1169 1417
rect 59 1398 1085 1404
rect 0 1386 1085 1398
rect 0 1334 7 1386
rect 59 1376 1085 1386
rect 59 1334 66 1376
rect 1113 1353 1115 1405
rect 1167 1353 1169 1405
rect 2216 1404 2223 1450
rect 1197 1398 2223 1404
rect 2275 1398 2282 1450
rect 1197 1386 2282 1398
rect 1197 1376 2223 1386
rect 1113 1348 1169 1353
rect 0 1322 66 1334
rect 0 1270 7 1322
rect 59 1292 66 1322
rect 94 1341 2188 1348
rect 94 1320 1115 1341
rect 59 1270 1085 1292
rect 0 1225 1085 1270
rect 1113 1289 1115 1320
rect 1167 1320 2188 1341
rect 2216 1334 2223 1376
rect 2275 1334 2282 1386
rect 2216 1322 2282 1334
rect 1167 1289 1169 1320
rect 2216 1292 2223 1322
rect 1113 1277 1169 1289
rect 1113 1225 1115 1277
rect 1167 1225 1169 1277
rect 1197 1270 2223 1292
rect 2275 1270 2282 1322
rect 1197 1225 2282 1270
rect 0 1224 66 1225
rect 1113 1197 1169 1225
rect 2216 1224 2282 1225
rect 74 1196 2208 1197
rect 0 1195 2282 1196
rect 0 1143 152 1195
rect 204 1143 216 1195
rect 268 1143 280 1195
rect 332 1143 344 1195
rect 396 1143 408 1195
rect 460 1143 472 1195
rect 524 1143 536 1195
rect 588 1143 600 1195
rect 652 1143 664 1195
rect 716 1143 728 1195
rect 780 1143 792 1195
rect 844 1143 856 1195
rect 908 1143 920 1195
rect 972 1143 984 1195
rect 1036 1143 1048 1195
rect 1100 1143 1182 1195
rect 1234 1143 1246 1195
rect 1298 1143 1310 1195
rect 1362 1143 1374 1195
rect 1426 1143 1438 1195
rect 1490 1143 1502 1195
rect 1554 1143 1566 1195
rect 1618 1143 1630 1195
rect 1682 1143 1694 1195
rect 1746 1143 1758 1195
rect 1810 1143 1822 1195
rect 1874 1143 1886 1195
rect 1938 1143 1950 1195
rect 2002 1143 2014 1195
rect 2066 1143 2078 1195
rect 2130 1143 2282 1195
rect 0 1142 2282 1143
rect 74 1141 2208 1142
rect 0 1113 66 1114
rect 1113 1113 1169 1141
rect 2216 1113 2282 1114
rect 0 1068 1085 1113
rect 0 1016 7 1068
rect 59 1046 1085 1068
rect 1113 1061 1115 1113
rect 1167 1061 1169 1113
rect 1113 1049 1169 1061
rect 59 1016 66 1046
rect 1113 1018 1115 1049
rect 0 1004 66 1016
rect 0 952 7 1004
rect 59 962 66 1004
rect 94 997 1115 1018
rect 1167 1018 1169 1049
rect 1197 1068 2282 1113
rect 1197 1046 2223 1068
rect 1167 997 2188 1018
rect 94 990 2188 997
rect 2216 1016 2223 1046
rect 2275 1016 2282 1068
rect 2216 1004 2282 1016
rect 1113 985 1169 990
rect 59 952 1085 962
rect 0 940 1085 952
rect 0 888 7 940
rect 59 934 1085 940
rect 59 888 66 934
rect 1113 933 1115 985
rect 1167 933 1169 985
rect 2216 962 2223 1004
rect 1197 952 2223 962
rect 2275 952 2282 1004
rect 1197 940 2282 952
rect 1197 934 2223 940
rect 1113 921 1169 933
rect 1113 906 1115 921
rect 0 876 66 888
rect 94 878 1115 906
rect 0 824 7 876
rect 59 850 66 876
rect 1113 869 1115 878
rect 1167 906 1169 921
rect 1167 878 2188 906
rect 2216 888 2223 934
rect 2275 888 2282 940
rect 1167 869 1169 878
rect 1113 857 1169 869
rect 59 824 1085 850
rect 0 822 1085 824
rect 0 812 66 822
rect 0 760 7 812
rect 59 760 66 812
rect 1113 805 1115 857
rect 1167 805 1169 857
rect 2216 876 2282 888
rect 2216 850 2223 876
rect 1197 824 2223 850
rect 2275 824 2282 876
rect 1197 822 2282 824
rect 1113 794 1169 805
rect 2216 812 2282 822
rect 94 793 2188 794
rect 94 766 1115 793
rect 0 748 66 760
rect 0 696 7 748
rect 59 738 66 748
rect 1113 741 1115 766
rect 1167 766 2188 793
rect 1167 741 1169 766
rect 59 710 1085 738
rect 1113 729 1169 741
rect 2216 760 2223 812
rect 2275 760 2282 812
rect 2216 748 2282 760
rect 2216 738 2223 748
rect 59 696 66 710
rect 0 684 66 696
rect 0 632 7 684
rect 59 632 66 684
rect 1113 682 1115 729
rect 94 677 1115 682
rect 1167 682 1169 729
rect 1197 710 2223 738
rect 2216 696 2223 710
rect 2275 696 2282 748
rect 2216 684 2282 696
rect 1167 677 2188 682
rect 94 665 2188 677
rect 94 654 1115 665
rect 0 626 66 632
rect 0 620 1085 626
rect 0 568 7 620
rect 59 598 1085 620
rect 1113 613 1115 654
rect 1167 654 2188 665
rect 1167 613 1169 654
rect 2216 632 2223 684
rect 2275 632 2282 684
rect 2216 626 2282 632
rect 1113 601 1169 613
rect 59 568 66 598
rect 1113 570 1115 601
rect 0 556 66 568
rect 0 504 7 556
rect 59 514 66 556
rect 94 549 1115 570
rect 1167 570 1169 601
rect 1197 620 2282 626
rect 1197 598 2223 620
rect 1167 549 2188 570
rect 94 542 2188 549
rect 2216 568 2223 598
rect 2275 568 2282 620
rect 2216 556 2282 568
rect 1113 537 1169 542
rect 59 504 1085 514
rect 0 492 1085 504
rect 0 440 7 492
rect 59 486 1085 492
rect 59 440 66 486
rect 1113 485 1115 537
rect 1167 485 1169 537
rect 2216 514 2223 556
rect 1197 504 2223 514
rect 2275 504 2282 556
rect 1197 492 2282 504
rect 1197 486 2223 492
rect 1113 473 1169 485
rect 1113 458 1115 473
rect 0 428 66 440
rect 94 430 1115 458
rect 0 376 7 428
rect 59 402 66 428
rect 1113 421 1115 430
rect 1167 458 1169 473
rect 1167 430 2188 458
rect 2216 440 2223 486
rect 2275 440 2282 492
rect 1167 421 1169 430
rect 1113 409 1169 421
rect 59 376 1085 402
rect 0 374 1085 376
rect 0 364 66 374
rect 0 312 7 364
rect 59 312 66 364
rect 1113 357 1115 409
rect 1167 357 1169 409
rect 2216 428 2282 440
rect 2216 402 2223 428
rect 1197 376 2223 402
rect 2275 376 2282 428
rect 1197 374 2282 376
rect 1113 346 1169 357
rect 2216 364 2282 374
rect 94 345 2188 346
rect 94 318 1115 345
rect 0 300 66 312
rect 0 248 7 300
rect 59 290 66 300
rect 1113 293 1115 318
rect 1167 318 2188 345
rect 1167 293 1169 318
rect 59 262 1085 290
rect 1113 281 1169 293
rect 2216 312 2223 364
rect 2275 312 2282 364
rect 2216 300 2282 312
rect 2216 290 2223 300
rect 59 248 66 262
rect 0 236 66 248
rect 0 184 7 236
rect 59 184 66 236
rect 1113 234 1115 281
rect 94 229 1115 234
rect 1167 234 1169 281
rect 1197 262 2223 290
rect 2216 248 2223 262
rect 2275 248 2282 300
rect 2216 236 2282 248
rect 1167 229 2188 234
rect 94 217 2188 229
rect 94 206 1115 217
rect 0 178 66 184
rect 0 172 1085 178
rect 0 120 7 172
rect 59 150 1085 172
rect 1113 165 1115 206
rect 1167 206 2188 217
rect 1167 165 1169 206
rect 2216 184 2223 236
rect 2275 184 2282 236
rect 2216 178 2282 184
rect 1113 153 1169 165
rect 59 120 66 150
rect 1113 122 1115 153
rect 0 108 66 120
rect 0 56 7 108
rect 59 66 66 108
rect 94 101 1115 122
rect 1167 122 1169 153
rect 1197 172 2282 178
rect 1197 150 2223 172
rect 1167 101 2188 122
rect 94 94 2188 101
rect 2216 120 2223 150
rect 2275 120 2282 172
rect 2216 108 2282 120
rect 59 59 1086 66
rect 59 56 88 59
rect 0 7 88 56
rect 140 7 152 59
rect 204 7 216 59
rect 268 7 280 59
rect 332 7 344 59
rect 396 7 408 59
rect 460 7 472 59
rect 524 7 536 59
rect 588 7 600 59
rect 652 7 664 59
rect 716 7 728 59
rect 780 7 792 59
rect 844 7 856 59
rect 908 7 920 59
rect 972 7 984 59
rect 1036 7 1086 59
rect 0 0 1086 7
rect 1114 0 1168 94
rect 2216 66 2223 108
rect 1196 59 2223 66
rect 1196 7 1246 59
rect 1298 7 1310 59
rect 1362 7 1374 59
rect 1426 7 1438 59
rect 1490 7 1502 59
rect 1554 7 1566 59
rect 1618 7 1630 59
rect 1682 7 1694 59
rect 1746 7 1758 59
rect 1810 7 1822 59
rect 1874 7 1886 59
rect 1938 7 1950 59
rect 2002 7 2014 59
rect 2066 7 2078 59
rect 2130 7 2142 59
rect 2194 56 2223 59
rect 2275 56 2282 108
rect 2194 7 2282 56
rect 1196 0 2282 7
<< labels >>
flabel metal2 s 1019 2162 1049 2184 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 1121 2062 1163 2098 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 1176 1289 1197 1338 0 FreeSans 1600 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 773906
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 748772
string gencell sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield
string library sky130
string parameter m=1
string device primitive
<< end >>
