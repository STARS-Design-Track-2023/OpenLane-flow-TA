magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 734 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 155 47 185 177
rect 351 47 381 177
rect 447 47 477 177
rect 540 47 570 177
rect 624 47 654 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 351 297 381 497
rect 447 297 477 497
rect 540 297 570 497
rect 624 297 654 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 47 155 177
rect 185 101 237 177
rect 185 67 195 101
rect 229 67 237 101
rect 185 47 237 67
rect 299 101 351 177
rect 299 67 307 101
rect 341 67 351 101
rect 299 47 351 67
rect 381 47 447 177
rect 477 97 540 177
rect 477 63 487 97
rect 521 63 540 97
rect 477 47 540 63
rect 570 101 624 177
rect 570 67 580 101
rect 614 67 624 101
rect 570 47 624 67
rect 654 165 708 177
rect 654 131 666 165
rect 700 131 708 165
rect 654 97 708 131
rect 654 63 666 97
rect 700 63 708 97
rect 654 47 708 63
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 409 163 497
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 485 245 497
rect 193 451 203 485
rect 237 451 245 485
rect 193 297 245 451
rect 299 477 351 497
rect 299 443 307 477
rect 341 443 351 477
rect 299 297 351 443
rect 381 477 447 497
rect 381 443 396 477
rect 430 443 447 477
rect 381 407 447 443
rect 381 373 396 407
rect 430 373 447 407
rect 381 297 447 373
rect 477 477 540 497
rect 477 443 496 477
rect 530 443 540 477
rect 477 409 540 443
rect 477 375 496 409
rect 530 375 540 409
rect 477 297 540 375
rect 570 477 624 497
rect 570 443 580 477
rect 614 443 624 477
rect 570 409 624 443
rect 570 375 580 409
rect 614 375 624 409
rect 570 297 624 375
rect 654 479 708 497
rect 654 445 666 479
rect 700 445 708 479
rect 654 411 708 445
rect 654 377 666 411
rect 700 377 708 411
rect 654 343 708 377
rect 654 309 666 343
rect 700 309 708 343
rect 654 297 708 309
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 195 67 229 101
rect 307 67 341 101
rect 487 63 521 97
rect 580 67 614 101
rect 666 131 700 165
rect 666 63 700 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 375 153 409
rect 203 451 237 485
rect 307 443 341 477
rect 396 443 430 477
rect 396 373 430 407
rect 496 443 530 477
rect 496 375 530 409
rect 580 443 614 477
rect 580 375 614 409
rect 666 445 700 479
rect 666 377 700 411
rect 666 309 700 343
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 351 497 381 523
rect 447 497 477 523
rect 540 497 570 523
rect 624 497 654 523
rect 79 265 109 297
rect 163 265 193 297
rect 351 265 381 297
rect 447 265 477 297
rect 540 265 570 297
rect 624 265 654 297
rect 55 249 109 265
rect 55 215 65 249
rect 99 215 109 249
rect 55 199 109 215
rect 79 177 109 199
rect 155 249 213 265
rect 155 215 169 249
rect 203 215 213 249
rect 155 199 213 215
rect 308 249 381 265
rect 308 215 318 249
rect 352 215 381 249
rect 308 199 381 215
rect 423 249 477 265
rect 423 215 433 249
rect 467 215 477 249
rect 423 199 477 215
rect 519 249 654 265
rect 519 215 529 249
rect 563 215 654 249
rect 519 199 654 215
rect 155 177 185 199
rect 351 177 381 199
rect 447 177 477 199
rect 540 177 570 199
rect 624 177 654 199
rect 79 21 109 47
rect 155 21 185 47
rect 351 21 381 47
rect 447 21 477 47
rect 540 21 570 47
rect 624 21 654 47
<< polycont >>
rect 65 215 99 249
rect 169 215 203 249
rect 318 215 352 249
rect 433 215 467 249
rect 529 215 563 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 19 485 253 493
rect 19 451 35 485
rect 69 459 203 485
rect 69 451 85 459
rect 187 451 203 459
rect 237 451 253 485
rect 291 477 362 527
rect 19 417 85 451
rect 291 443 307 477
rect 341 443 362 477
rect 396 477 446 493
rect 430 443 446 477
rect 19 383 35 417
rect 69 383 85 417
rect 19 349 85 383
rect 119 409 165 425
rect 153 407 165 409
rect 396 407 446 443
rect 153 375 396 407
rect 119 373 396 375
rect 430 373 446 407
rect 480 477 546 527
rect 480 443 496 477
rect 530 443 546 477
rect 480 409 546 443
rect 480 375 496 409
rect 530 375 546 409
rect 580 477 632 493
rect 614 443 632 477
rect 580 409 632 443
rect 614 375 632 409
rect 119 359 446 373
rect 580 357 632 375
rect 19 315 35 349
rect 69 325 85 349
rect 69 315 563 325
rect 19 291 563 315
rect 18 249 115 255
rect 18 215 65 249
rect 99 215 115 249
rect 153 249 248 257
rect 153 215 169 249
rect 203 215 248 249
rect 19 165 109 170
rect 19 131 35 165
rect 69 131 109 165
rect 204 135 248 215
rect 302 249 368 257
rect 302 215 318 249
rect 352 215 368 249
rect 402 249 483 255
rect 402 215 433 249
rect 467 215 483 249
rect 529 249 563 291
rect 302 135 344 215
rect 529 181 563 215
rect 395 147 563 181
rect 19 97 109 131
rect 395 101 429 147
rect 598 117 632 357
rect 666 479 700 527
rect 666 411 700 445
rect 666 343 700 377
rect 666 289 700 309
rect 19 63 35 97
rect 69 63 109 97
rect 19 17 109 63
rect 164 67 195 101
rect 229 67 307 101
rect 341 67 429 101
rect 164 51 429 67
rect 471 97 537 113
rect 471 63 487 97
rect 521 63 537 97
rect 471 17 537 63
rect 580 101 632 117
rect 614 67 632 101
rect 580 51 632 67
rect 666 165 700 197
rect 666 97 700 131
rect 666 17 700 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 310 221 344 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 402 221 436 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 586 425 620 459 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 310 153 344 187 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 214 153 248 187 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 586 357 620 391 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a22o_2
rlabel metal1 s 0 -48 736 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 4059210
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4052462
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 18.400 0.000 
<< end >>
