magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__dfl1sd2__example_5595914180812  sky130_fd_pr__dfl1sd2__example_5595914180812_0
timestamp 1686671242
transform 1 0 50 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180811  sky130_fd_pr__dfl1sd__example_5595914180811_0
timestamp 1686671242
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180811  sky130_fd_pr__dfl1sd__example_5595914180811_1
timestamp 1686671242
transform 1 0 156 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 6905982
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6904482
<< end >>
