magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -36 679 836 1471
<< pwell >>
rect 664 25 766 159
<< psubdiff >>
rect 690 109 740 133
rect 690 75 698 109
rect 732 75 740 109
rect 690 51 740 75
<< nsubdiff >>
rect 690 1339 740 1363
rect 690 1305 698 1339
rect 732 1305 740 1339
rect 690 1281 740 1305
<< psubdiffcont >>
rect 698 75 732 109
<< nsubdiffcont >>
rect 698 1305 732 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 800 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 698 1339 732 1397
rect 698 1289 732 1305
rect 64 724 98 740
rect 64 674 98 690
rect 380 724 414 1096
rect 380 690 431 724
rect 380 318 414 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 698 109 732 125
rect 698 17 732 75
rect 0 -17 800 17
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1686671242
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_28  sky130_sram_2kbyte_1rw1r_32x512_8_contact_28_0
timestamp 1686671242
transform 1 0 690 0 1 1281
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_29  sky130_sram_2kbyte_1rw1r_32x512_8_contact_29_0
timestamp 1686671242
transform 1 0 690 0 1 51
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m5_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m5_w2_000_sli_dli_da_p_0
timestamp 1686671242
transform 1 0 54 0 1 51
box -26 -26 608 456
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m5_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m5_w2_000_sli_dli_da_p_0
timestamp 1686671242
transform 1 0 54 0 1 963
box -59 -56 641 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 414 707 414 707 4 Z
rlabel locali s 400 0 400 0 4 gnd
rlabel locali s 400 1414 400 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 800 1414
string GDS_END 390336
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 388210
<< end >>
