magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< locali >>
rect 12028 18138 12590 18733
rect 1835 1730 2397 2325
rect 1835 -41064 2397 -40469
<< obsli1 >>
rect 12922 20881 13056 20947
rect 13222 20881 13356 20947
rect 12886 20781 12920 20847
rect 12972 20781 13006 20847
rect 13058 20781 13092 20847
rect 13186 20781 13220 20847
rect 13272 20781 13306 20847
rect 13358 20781 13392 20847
rect 14491 20240 14525 20810
rect 14577 20240 14611 20810
rect 14663 20240 14697 20810
rect 14749 20240 14783 20810
rect 14835 20240 14869 20810
rect 14921 20240 14955 20810
rect 15007 20240 15041 20810
rect 15093 20240 15127 20810
rect 15179 20240 15213 20810
rect 15307 20240 15341 20810
rect 15393 20240 15427 20810
rect 15479 20240 15513 20810
rect 15565 20240 15599 20810
rect 15651 20240 15685 20810
rect 15737 20240 15771 20810
rect 15823 20240 15857 20810
rect 15909 20240 15943 20810
rect 15995 20240 16029 20810
rect 20992 20767 21026 20905
rect 21078 20767 21112 20905
rect 21164 20767 21198 20905
rect 21250 20767 21284 20905
rect 21336 20767 21370 20905
rect 20099 20671 20133 20737
rect 20185 20671 20219 20737
rect 20271 20671 20305 20737
rect 21046 20655 21316 20721
rect 22641 20698 22675 21268
rect 22727 20698 22761 21268
rect 22813 20698 22847 21268
rect 22899 20698 22933 21268
rect 22985 20698 23019 21268
rect 23071 20698 23105 21268
rect 23157 20698 23191 21268
rect 23243 20698 23277 21268
rect 23329 20698 23363 21268
rect 19853 20571 19987 20637
rect 20135 20571 20269 20637
rect 19817 20471 19851 20537
rect 19903 20471 19937 20537
rect 19989 20471 20023 20537
rect 20099 20471 20133 20537
rect 20185 20471 20219 20537
rect 20271 20471 20305 20537
rect 20992 20471 21026 20609
rect 21078 20471 21112 20609
rect 21164 20471 21198 20609
rect 21250 20471 21284 20609
rect 21336 20471 21370 20609
rect 22731 20586 23273 20652
rect 22899 20486 22933 20552
rect 22985 20486 23019 20552
rect 23071 20486 23105 20552
rect 14581 20128 15123 20194
rect 15397 20128 15939 20194
rect 15362 -24034 15496 -23968
rect 15656 -24034 15790 -23968
rect 13728 -24867 13862 -24799
rect 14028 -24867 14162 -24799
rect 13692 -25051 13726 -24913
rect 13778 -25051 13812 -24913
rect 13864 -25051 13898 -24913
rect 13992 -25051 14026 -24913
rect 14078 -25051 14112 -24913
rect 14164 -25051 14198 -24913
rect 15326 -25066 15360 -24068
rect 15412 -25066 15446 -24068
rect 15498 -25066 15532 -24068
rect 15620 -25066 15654 -24068
rect 15706 -25066 15740 -24068
rect 15792 -25066 15826 -24068
rect 21549 -24583 21583 -24277
rect 21635 -24583 21669 -24277
rect 21721 -24583 21755 -24277
rect 21807 -24583 21841 -24277
rect 21893 -24583 21927 -24277
rect 23371 -24583 23405 -24277
rect 23457 -24583 23491 -24277
rect 23543 -24583 23577 -24277
rect 23629 -24583 23663 -24277
rect 23715 -24583 23749 -24277
rect 20186 -24751 20220 -24613
rect 20272 -24751 20306 -24613
rect 20358 -24751 20392 -24613
rect 21603 -24699 21873 -24629
rect 22051 -24699 22321 -24631
rect 23425 -24697 23695 -24629
rect 20222 -24867 20356 -24797
rect 20186 -25051 20220 -24913
rect 20272 -25051 20306 -24913
rect 20358 -25051 20392 -24913
rect 21549 -25051 21583 -24745
rect 21635 -25051 21669 -24745
rect 21721 -25051 21755 -24745
rect 21807 -25051 21841 -24745
rect 21893 -25051 21927 -24745
rect 21997 -25051 22031 -24745
rect 22083 -25051 22117 -24745
rect 22169 -25051 22203 -24745
rect 22255 -25051 22289 -24745
rect 22341 -25051 22375 -24745
rect 23457 -25729 23491 -24731
rect 23543 -25729 23577 -24731
rect 23629 -25729 23663 -24731
<< obsm1 >>
rect 22635 21348 23369 21408
rect 20986 20985 21376 21045
rect 12924 20885 13054 20943
rect 13224 20885 13354 20943
rect 14485 20890 15219 20950
rect 12880 20701 12926 20850
rect 12963 20781 13015 20850
rect 13052 20701 13098 20850
rect 12880 20641 13098 20701
rect 13180 20701 13226 20850
rect 13263 20781 13315 20850
rect 13352 20701 13398 20850
rect 13180 20641 13398 20701
rect 14485 20240 14531 20890
rect 14568 20240 14620 20810
rect 14657 20240 14703 20890
rect 14740 20240 14792 20810
rect 14829 20240 14875 20890
rect 14912 20240 14964 20810
rect 15001 20240 15047 20890
rect 15084 20240 15136 20810
rect 15173 20240 15219 20890
rect 15301 20890 16035 20950
rect 15301 20240 15347 20890
rect 15384 20240 15436 20810
rect 15473 20240 15519 20890
rect 15556 20240 15608 20810
rect 15645 20240 15691 20890
rect 15728 20240 15780 20810
rect 15817 20240 15863 20890
rect 15900 20240 15952 20810
rect 15989 20240 16035 20890
rect 20093 20817 20311 20877
rect 20093 20668 20139 20817
rect 20176 20668 20228 20737
rect 20265 20668 20311 20817
rect 20986 20767 21032 20985
rect 21069 20767 21121 20905
rect 21158 20767 21204 20985
rect 21241 20767 21293 20905
rect 21330 20767 21376 20985
rect 21044 20659 21318 20717
rect 22635 20698 22681 21348
rect 22718 20698 22770 21268
rect 22807 20698 22853 21348
rect 22890 20698 22942 21268
rect 22979 20698 23025 21348
rect 23062 20698 23114 21268
rect 23151 20698 23197 21348
rect 23234 20698 23286 21268
rect 23323 20698 23369 21348
rect 19855 20575 19985 20633
rect 20137 20575 20267 20633
rect 19811 20391 19857 20540
rect 19894 20471 19946 20540
rect 19983 20391 20029 20540
rect 19811 20331 20029 20391
rect 20093 20391 20139 20540
rect 20176 20471 20228 20540
rect 20265 20391 20311 20540
rect 20093 20331 20311 20391
rect 20986 20391 21032 20609
rect 21069 20471 21121 20609
rect 21158 20391 21204 20609
rect 21241 20471 21293 20609
rect 21330 20391 21376 20609
rect 22721 20590 23283 20648
rect 20986 20331 21376 20391
rect 22893 20406 22939 20555
rect 22976 20486 23028 20555
rect 23065 20406 23111 20555
rect 22893 20346 23111 20406
rect 14571 20132 15133 20190
rect 15387 20132 15949 20190
rect 15364 -24030 15494 -23972
rect 15658 -24030 15788 -23972
rect 13730 -24861 13860 -24803
rect 14030 -24861 14160 -24803
rect 13686 -25131 13732 -24913
rect 13769 -25051 13821 -24913
rect 13858 -25131 13904 -24913
rect 13686 -25191 13904 -25131
rect 13986 -25131 14032 -24913
rect 14069 -25051 14121 -24913
rect 14158 -25131 14204 -24913
rect 13986 -25191 14204 -25131
rect 15320 -25147 15366 -24068
rect 15403 -25066 15455 -24068
rect 15492 -25147 15538 -24068
rect 15320 -25199 15538 -25147
rect 15614 -25147 15660 -24068
rect 15697 -25066 15749 -24068
rect 15786 -25147 15832 -24068
rect 21543 -24197 21933 -24137
rect 20180 -24533 20398 -24473
rect 20180 -24751 20226 -24533
rect 20263 -24751 20315 -24613
rect 20352 -24751 20398 -24533
rect 21543 -24583 21589 -24197
rect 21626 -24583 21678 -24277
rect 21715 -24583 21761 -24197
rect 21798 -24583 21850 -24277
rect 21887 -24583 21933 -24197
rect 23365 -24197 23755 -24137
rect 23365 -24583 23411 -24197
rect 23448 -24583 23500 -24277
rect 23537 -24583 23583 -24197
rect 23620 -24583 23672 -24277
rect 23709 -24583 23755 -24197
rect 21601 -24693 21875 -24635
rect 22049 -24693 22323 -24635
rect 23423 -24693 23697 -24635
rect 20224 -24861 20354 -24803
rect 15614 -25199 15832 -25147
rect 20180 -25131 20226 -24913
rect 20263 -25051 20315 -24913
rect 20352 -25131 20398 -24913
rect 20180 -25191 20398 -25131
rect 21543 -25131 21589 -24745
rect 21626 -25051 21678 -24745
rect 21715 -25131 21761 -24745
rect 21798 -25051 21850 -24745
rect 21887 -25131 21933 -24745
rect 21543 -25191 21933 -25131
rect 21991 -25131 22037 -24745
rect 22074 -25051 22126 -24745
rect 22163 -25131 22209 -24745
rect 22246 -25051 22298 -24745
rect 22335 -25131 22381 -24745
rect 21991 -25191 22381 -25131
rect 23451 -25810 23497 -24731
rect 23534 -25729 23586 -24731
rect 23623 -25810 23669 -24731
rect 23451 -25862 23669 -25810
<< obsm2 >>
rect 12963 20781 13015 20850
rect 13263 20781 13315 20850
rect 21062 20761 21128 20915
rect 21234 20761 21300 20915
rect 20176 20668 20228 20737
rect 22711 20692 22777 20846
rect 22883 20692 22949 20846
rect 23055 20692 23121 20846
rect 23227 20692 23293 20846
rect 19894 20471 19946 20540
rect 20176 20471 20228 20540
rect 21062 20461 21128 20615
rect 21234 20461 21300 20615
rect 22976 20486 23028 20555
rect 14561 20234 14627 20388
rect 14733 20234 14799 20388
rect 14905 20234 14971 20388
rect 15077 20234 15143 20388
rect 15377 20234 15443 20388
rect 15549 20234 15615 20388
rect 15721 20234 15787 20388
rect 15893 20234 15959 20388
rect 15403 -24198 15455 -24070
rect 15697 -24198 15749 -24070
rect 21619 -24591 21685 -24437
rect 21791 -24591 21857 -24437
rect 23441 -24591 23507 -24437
rect 23613 -24591 23679 -24437
rect 20263 -24746 20315 -24618
rect 21619 -24891 21685 -24737
rect 21791 -24891 21857 -24737
rect 22067 -24891 22133 -24737
rect 22239 -24891 22305 -24737
rect 23534 -24861 23586 -24733
rect 13769 -25046 13821 -24918
rect 14069 -25046 14121 -24918
rect 20263 -25046 20315 -24918
<< obsm3 >>
rect 21062 20827 21128 20915
rect 21234 20827 21300 20915
rect 21062 20761 21300 20827
rect 22711 20758 22777 20846
rect 22883 20758 22949 20846
rect 23055 20758 23121 20846
rect 23227 20758 23293 20846
rect 22711 20692 23293 20758
rect 21062 20549 21300 20615
rect 21062 20461 21128 20549
rect 21234 20461 21300 20549
rect 14561 20300 14627 20388
rect 14733 20300 14799 20388
rect 14905 20300 14971 20388
rect 15077 20300 15143 20388
rect 14561 20234 15143 20300
rect 15377 20300 15443 20388
rect 15549 20300 15615 20388
rect 15721 20300 15787 20388
rect 15893 20300 15959 20388
rect 15377 20234 15959 20300
rect 21619 -24525 21685 -24437
rect 21791 -24525 21857 -24437
rect 21619 -24591 21857 -24525
rect 23441 -24525 23507 -24437
rect 23613 -24525 23679 -24437
rect 23441 -24591 23679 -24525
rect 21619 -24803 21857 -24737
rect 21619 -24891 21685 -24803
rect 21791 -24891 21857 -24803
rect 22067 -24803 22305 -24737
rect 22067 -24891 22133 -24803
rect 22239 -24891 22305 -24803
<< labels >>
rlabel locali s 1835 -41064 2397 -40469 8 B_P
port 1 nsew
rlabel locali s 1835 1730 2397 2325 6 NWELL
port 2 nsew
rlabel locali s 12028 18138 12590 18733 6 VGND
port 3 nsew ground default
<< properties >>
string FIXED_BBOX 0 -42794 311106 39640
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10508798
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10504344
<< end >>
