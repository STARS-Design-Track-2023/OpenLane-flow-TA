magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -36 679 294 1471
<< poly >>
rect 114 740 144 937
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 477 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 258 1431
rect 62 1130 96 1397
rect 64 724 98 740
rect 64 674 98 690
rect 162 724 196 1196
rect 162 690 213 724
rect 162 218 196 690
rect 62 17 96 218
rect 0 -17 258 17
use contact_12  contact_12_0
timestamp 1686671242
transform 1 0 48 0 1 674
box 0 0 1 1
use nmos_m13_w2_000_sli_dli_da_p  nmos_m13_w2_000_sli_dli_da_p_0
timestamp 1686671242
transform 1 0 54 0 1 51
box -26 -26 176 426
use pmos_m13_w2_000_sli_dli_da_p  pmos_m13_w2_000_sli_dli_da_p_0
timestamp 1686671242
transform 1 0 54 0 1 963
box -59 -54 209 454
<< labels >>
rlabel locali s 196 707 196 707 4 Z
port 2 nsew
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 129 1414 129 1414 4 vdd
port 3 nsew
rlabel locali s 129 0 129 0 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 258 1414
string GDS_END 3373780
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 3372386
<< end >>
