magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__dfm1sd2__example_55959141808219  sky130_fd_pr__dfm1sd2__example_55959141808219_0
timestamp 1686671242
transform 1 0 200 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd__example_55959141808225  sky130_fd_pr__dfm1sd__example_55959141808225_0
timestamp 1686671242
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808207  sky130_fd_pr__hvdfm1sd__example_55959141808207_0
timestamp 1686671242
transform 1 0 456 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 37270168
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37268728
<< end >>
