magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 133 157 919 203
rect 36 21 919 157
rect 36 17 58 21
rect 24 -17 58 17
<< locali >>
rect 17 199 114 340
rect 532 335 621 493
rect 532 299 713 335
rect 547 199 713 299
rect 547 165 621 199
rect 532 51 621 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 408 104 493
rect 138 442 215 527
rect 17 374 215 408
rect 148 265 215 374
rect 249 335 303 493
rect 337 408 387 493
rect 421 442 498 527
rect 337 369 498 408
rect 249 299 394 335
rect 148 199 230 265
rect 264 199 394 299
rect 428 265 498 369
rect 655 408 706 493
rect 740 442 817 527
rect 655 369 817 408
rect 428 199 513 265
rect 747 265 817 369
rect 851 299 903 493
rect 747 199 832 265
rect 148 165 215 199
rect 264 165 303 199
rect 428 165 498 199
rect 747 165 817 199
rect 866 165 903 299
rect 17 131 215 165
rect 17 51 104 131
rect 138 17 215 97
rect 249 51 303 165
rect 337 131 498 165
rect 337 51 387 131
rect 421 17 498 97
rect 655 131 817 165
rect 655 51 706 131
rect 740 17 817 97
rect 851 51 903 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 17 199 114 340 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 920 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 24 -17 58 17 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 36 17 58 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 36 21 919 157 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 133 157 919 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 532 51 621 165 6 X
port 6 nsew signal output
rlabel locali s 547 165 621 199 6 X
port 6 nsew signal output
rlabel locali s 547 199 713 299 6 X
port 6 nsew signal output
rlabel locali s 532 299 713 335 6 X
port 6 nsew signal output
rlabel locali s 532 335 621 493 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 920 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2925094
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2917318
<< end >>
