magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< pwell >>
rect 10 76 686 458
<< nmos >>
rect 204 102 234 432
rect 290 102 320 432
rect 376 102 406 432
rect 462 102 492 432
<< ndiff >>
rect 148 420 204 432
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 234 420 290 432
rect 234 386 245 420
rect 279 386 290 420
rect 234 352 290 386
rect 234 318 245 352
rect 279 318 290 352
rect 234 284 290 318
rect 234 250 245 284
rect 279 250 290 284
rect 234 216 290 250
rect 234 182 245 216
rect 279 182 290 216
rect 234 148 290 182
rect 234 114 245 148
rect 279 114 290 148
rect 234 102 290 114
rect 320 420 376 432
rect 320 386 331 420
rect 365 386 376 420
rect 320 352 376 386
rect 320 318 331 352
rect 365 318 376 352
rect 320 284 376 318
rect 320 250 331 284
rect 365 250 376 284
rect 320 216 376 250
rect 320 182 331 216
rect 365 182 376 216
rect 320 148 376 182
rect 320 114 331 148
rect 365 114 376 148
rect 320 102 376 114
rect 406 420 462 432
rect 406 386 417 420
rect 451 386 462 420
rect 406 352 462 386
rect 406 318 417 352
rect 451 318 462 352
rect 406 284 462 318
rect 406 250 417 284
rect 451 250 462 284
rect 406 216 462 250
rect 406 182 417 216
rect 451 182 462 216
rect 406 148 462 182
rect 406 114 417 148
rect 451 114 462 148
rect 406 102 462 114
rect 492 420 548 432
rect 492 386 503 420
rect 537 386 548 420
rect 492 352 548 386
rect 492 318 503 352
rect 537 318 548 352
rect 492 284 548 318
rect 492 250 503 284
rect 537 250 548 284
rect 492 216 548 250
rect 492 182 503 216
rect 537 182 548 216
rect 492 148 548 182
rect 492 114 503 148
rect 537 114 548 148
rect 492 102 548 114
<< ndiffc >>
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 245 386 279 420
rect 245 318 279 352
rect 245 250 279 284
rect 245 182 279 216
rect 245 114 279 148
rect 331 386 365 420
rect 331 318 365 352
rect 331 250 365 284
rect 331 182 365 216
rect 331 114 365 148
rect 417 386 451 420
rect 417 318 451 352
rect 417 250 451 284
rect 417 182 451 216
rect 417 114 451 148
rect 503 386 537 420
rect 503 318 537 352
rect 503 250 537 284
rect 503 182 537 216
rect 503 114 537 148
<< psubdiff >>
rect 36 386 94 432
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 602 386 660 432
rect 602 352 614 386
rect 648 352 660 386
rect 602 318 660 352
rect 602 284 614 318
rect 648 284 660 318
rect 602 250 660 284
rect 602 216 614 250
rect 648 216 660 250
rect 602 182 660 216
rect 602 148 614 182
rect 648 148 660 182
rect 602 102 660 148
<< psubdiffcont >>
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 614 352 648 386
rect 614 284 648 318
rect 614 216 648 250
rect 614 148 648 182
<< poly >>
rect 179 504 517 524
rect 179 470 195 504
rect 229 470 263 504
rect 297 470 331 504
rect 365 470 399 504
rect 433 470 467 504
rect 501 470 517 504
rect 179 454 517 470
rect 204 432 234 454
rect 290 432 320 454
rect 376 432 406 454
rect 462 432 492 454
rect 204 80 234 102
rect 290 80 320 102
rect 376 80 406 102
rect 462 80 492 102
rect 179 64 517 80
rect 179 30 195 64
rect 229 30 263 64
rect 297 30 331 64
rect 365 30 399 64
rect 433 30 467 64
rect 501 30 517 64
rect 179 10 517 30
<< polycont >>
rect 195 470 229 504
rect 263 470 297 504
rect 331 470 365 504
rect 399 470 433 504
rect 467 470 501 504
rect 195 30 229 64
rect 263 30 297 64
rect 331 30 365 64
rect 399 30 433 64
rect 467 30 501 64
<< locali >>
rect 179 470 187 504
rect 229 470 259 504
rect 297 470 331 504
rect 365 470 399 504
rect 437 470 467 504
rect 509 470 517 504
rect 159 420 193 436
rect 48 392 82 402
rect 48 320 82 352
rect 48 250 82 284
rect 48 182 82 214
rect 48 132 82 142
rect 159 352 193 358
rect 159 284 193 286
rect 159 248 193 250
rect 159 176 193 182
rect 159 98 193 114
rect 245 420 279 436
rect 245 352 279 358
rect 245 284 279 286
rect 245 248 279 250
rect 245 176 279 182
rect 245 98 279 114
rect 331 420 365 436
rect 331 352 365 358
rect 331 284 365 286
rect 331 248 365 250
rect 331 176 365 182
rect 331 98 365 114
rect 417 420 451 436
rect 417 352 451 358
rect 417 284 451 286
rect 417 248 451 250
rect 417 176 451 182
rect 417 98 451 114
rect 503 420 537 436
rect 503 352 537 358
rect 503 284 537 286
rect 503 248 537 250
rect 503 176 537 182
rect 614 392 648 402
rect 614 320 648 352
rect 614 250 648 284
rect 614 182 648 214
rect 614 132 648 142
rect 503 98 537 114
rect 179 30 187 64
rect 229 30 259 64
rect 297 30 331 64
rect 365 30 399 64
rect 437 30 467 64
rect 509 30 517 64
<< viali >>
rect 187 470 195 504
rect 195 470 221 504
rect 259 470 263 504
rect 263 470 293 504
rect 331 470 365 504
rect 403 470 433 504
rect 433 470 437 504
rect 475 470 501 504
rect 501 470 509 504
rect 48 386 82 392
rect 48 358 82 386
rect 48 318 82 320
rect 48 286 82 318
rect 48 216 82 248
rect 48 214 82 216
rect 48 148 82 176
rect 48 142 82 148
rect 159 386 193 392
rect 159 358 193 386
rect 159 318 193 320
rect 159 286 193 318
rect 159 216 193 248
rect 159 214 193 216
rect 159 148 193 176
rect 159 142 193 148
rect 245 386 279 392
rect 245 358 279 386
rect 245 318 279 320
rect 245 286 279 318
rect 245 216 279 248
rect 245 214 279 216
rect 245 148 279 176
rect 245 142 279 148
rect 331 386 365 392
rect 331 358 365 386
rect 331 318 365 320
rect 331 286 365 318
rect 331 216 365 248
rect 331 214 365 216
rect 331 148 365 176
rect 331 142 365 148
rect 417 386 451 392
rect 417 358 451 386
rect 417 318 451 320
rect 417 286 451 318
rect 417 216 451 248
rect 417 214 451 216
rect 417 148 451 176
rect 417 142 451 148
rect 503 386 537 392
rect 503 358 537 386
rect 503 318 537 320
rect 503 286 537 318
rect 503 216 537 248
rect 503 214 537 216
rect 503 148 537 176
rect 503 142 537 148
rect 614 386 648 392
rect 614 358 648 386
rect 614 318 648 320
rect 614 286 648 318
rect 614 216 648 248
rect 614 214 648 216
rect 614 148 648 176
rect 614 142 648 148
rect 187 30 195 64
rect 195 30 221 64
rect 259 30 263 64
rect 263 30 293 64
rect 331 30 365 64
rect 403 30 433 64
rect 433 30 437 64
rect 475 30 501 64
rect 501 30 509 64
<< metal1 >>
rect 175 504 521 524
rect 175 470 187 504
rect 221 470 259 504
rect 293 470 331 504
rect 365 470 403 504
rect 437 470 475 504
rect 509 470 521 504
rect 175 458 521 470
rect 36 392 94 420
rect 36 358 48 392
rect 82 358 94 392
rect 36 320 94 358
rect 36 286 48 320
rect 82 286 94 320
rect 36 248 94 286
rect 36 214 48 248
rect 82 214 94 248
rect 36 176 94 214
rect 36 142 48 176
rect 82 142 94 176
rect 36 114 94 142
rect 150 392 202 420
rect 150 358 159 392
rect 193 358 202 392
rect 150 320 202 358
rect 150 286 159 320
rect 193 286 202 320
rect 150 248 202 286
rect 150 236 159 248
rect 193 236 202 248
rect 150 176 202 184
rect 150 172 159 176
rect 193 172 202 176
rect 150 114 202 120
rect 236 414 288 420
rect 236 358 245 362
rect 279 358 288 362
rect 236 350 288 358
rect 236 286 245 298
rect 279 286 288 298
rect 236 248 288 286
rect 236 214 245 248
rect 279 214 288 248
rect 236 176 288 214
rect 236 142 245 176
rect 279 142 288 176
rect 236 114 288 142
rect 322 392 374 420
rect 322 358 331 392
rect 365 358 374 392
rect 322 320 374 358
rect 322 286 331 320
rect 365 286 374 320
rect 322 248 374 286
rect 322 236 331 248
rect 365 236 374 248
rect 322 176 374 184
rect 322 172 331 176
rect 365 172 374 176
rect 322 114 374 120
rect 408 414 460 420
rect 408 358 417 362
rect 451 358 460 362
rect 408 350 460 358
rect 408 286 417 298
rect 451 286 460 298
rect 408 248 460 286
rect 408 214 417 248
rect 451 214 460 248
rect 408 176 460 214
rect 408 142 417 176
rect 451 142 460 176
rect 408 114 460 142
rect 494 392 546 420
rect 494 358 503 392
rect 537 358 546 392
rect 494 320 546 358
rect 494 286 503 320
rect 537 286 546 320
rect 494 248 546 286
rect 494 236 503 248
rect 537 236 546 248
rect 494 176 546 184
rect 494 172 503 176
rect 537 172 546 176
rect 494 114 546 120
rect 602 392 660 420
rect 602 358 614 392
rect 648 358 660 392
rect 602 320 660 358
rect 602 286 614 320
rect 648 286 660 320
rect 602 248 660 286
rect 602 214 614 248
rect 648 214 660 248
rect 602 176 660 214
rect 602 142 614 176
rect 648 142 660 176
rect 602 114 660 142
rect 175 64 521 76
rect 175 30 187 64
rect 221 30 259 64
rect 293 30 331 64
rect 365 30 403 64
rect 437 30 475 64
rect 509 30 521 64
rect 175 10 521 30
<< via1 >>
rect 150 214 159 236
rect 159 214 193 236
rect 193 214 202 236
rect 150 184 202 214
rect 150 142 159 172
rect 159 142 193 172
rect 193 142 202 172
rect 150 120 202 142
rect 236 392 288 414
rect 236 362 245 392
rect 245 362 279 392
rect 279 362 288 392
rect 236 320 288 350
rect 236 298 245 320
rect 245 298 279 320
rect 279 298 288 320
rect 322 214 331 236
rect 331 214 365 236
rect 365 214 374 236
rect 322 184 374 214
rect 322 142 331 172
rect 331 142 365 172
rect 365 142 374 172
rect 322 120 374 142
rect 408 392 460 414
rect 408 362 417 392
rect 417 362 451 392
rect 451 362 460 392
rect 408 320 460 350
rect 408 298 417 320
rect 417 298 451 320
rect 451 298 460 320
rect 494 214 503 236
rect 503 214 537 236
rect 537 214 546 236
rect 494 184 546 214
rect 494 142 503 172
rect 503 142 537 172
rect 537 142 546 172
rect 494 120 546 142
<< metal2 >>
rect 10 414 686 420
rect 10 362 236 414
rect 288 362 408 414
rect 460 362 686 414
rect 10 350 686 362
rect 10 298 236 350
rect 288 298 408 350
rect 460 298 686 350
rect 10 292 686 298
rect 10 236 686 242
rect 10 184 150 236
rect 202 184 322 236
rect 374 184 494 236
rect 546 184 686 236
rect 10 172 686 184
rect 10 120 150 172
rect 202 120 322 172
rect 374 120 494 172
rect 546 120 686 172
rect 10 114 686 120
<< labels >>
flabel metal2 s 10 292 30 420 7 FreeSans 300 180 0 0 DRAIN
port 2 nsew
flabel metal2 s 10 114 30 242 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal1 s 602 114 660 130 3 FreeSans 300 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 175 458 521 524 0 FreeSans 300 0 0 0 GATE
port 5 nsew
flabel metal1 s 175 10 521 76 0 FreeSans 300 0 0 0 GATE
port 5 nsew
flabel metal1 s 36 114 94 130 3 FreeSans 300 90 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_END 5005564
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 4995168
<< end >>
