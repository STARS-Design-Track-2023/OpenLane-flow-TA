magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< metal4 >>
rect 0 35157 254 40000
rect 15746 35157 16000 40000
rect 0 14007 254 19000
rect 15746 14007 16000 19000
rect 0 12817 254 13707
rect 15746 12817 16000 13707
rect 0 11647 254 12537
rect 15746 11647 16000 12537
rect 0 11281 16000 11347
rect 0 10625 16000 11221
rect 0 10329 254 10565
rect 15746 10329 16000 10565
rect 0 9673 16000 10269
rect 0 9547 16000 9613
rect 0 8317 254 9247
rect 15746 8317 16000 9247
rect 0 7347 254 8037
rect 15746 7347 16000 8037
rect 0 6377 254 7067
rect 15746 6377 16000 7067
rect 0 5167 254 6097
rect 15746 5167 16000 6097
rect 0 3957 254 4887
rect 15746 3957 16000 4887
rect 0 2987 193 3677
rect 15794 2987 16000 3677
rect 0 1777 254 2707
rect 15746 1777 16000 2707
rect 0 407 254 1497
rect 15746 407 16000 1497
<< obsm4 >>
rect 334 35077 15666 40000
rect 193 19080 15794 35077
rect 334 13927 15666 19080
rect 193 13787 15794 13927
rect 334 12737 15666 13787
rect 193 12617 15794 12737
rect 334 11567 15666 12617
rect 193 11427 15794 11567
rect 334 10349 15666 10545
rect 193 9327 15794 9467
rect 334 8237 15666 9327
rect 193 8117 15794 8237
rect 334 7267 15666 8117
rect 193 7147 15794 7267
rect 334 6297 15666 7147
rect 193 6177 15794 6297
rect 334 5087 15666 6177
rect 193 4967 15794 5087
rect 334 3877 15666 4967
rect 193 3757 15794 3877
rect 273 2907 15714 3757
rect 193 2787 15794 2907
rect 334 1697 15666 2787
rect 193 1577 15794 1697
rect 334 407 15666 1577
<< metal5 >>
rect 0 35157 254 40000
rect 15746 35157 16000 40000
rect 2240 20912 14760 33392
rect 0 14007 254 18997
rect 0 12837 254 13687
rect 0 11667 254 12517
rect 0 9547 254 11347
rect 0 8337 254 9227
rect 0 7368 254 8017
rect 15746 14007 16000 18997
rect 15746 12837 16000 13687
rect 15746 11667 16000 12517
rect 15746 9547 16000 11347
rect 15746 8337 16000 9227
rect 15746 7368 16000 8017
rect 0 6397 254 7047
rect 0 5187 254 6077
rect 0 3977 254 4867
rect 15746 6397 16000 7047
rect 15746 5187 16000 6077
rect 15746 3977 16000 4867
rect 0 3007 193 3657
rect 15794 3007 16000 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 15746 1797 16000 2687
rect 15746 427 16000 1477
<< obsm5 >>
rect 574 34837 15426 40000
rect 0 33712 16000 34837
rect 0 20592 1920 33712
rect 15080 20592 16000 33712
rect 0 19317 16000 20592
rect 574 7368 15426 19317
rect 0 7367 16000 7368
rect 574 3657 15426 7367
rect 513 3007 15474 3657
rect 574 427 15426 3007
<< labels >>
rlabel metal5 s 2240 20912 14760 33392 6 PAD
port 1 nsew signal default
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 2 nsew ground bidirectional
rlabel metal5 s 15746 35157 16000 40000 6 VSSIO
port 2 nsew ground bidirectional
rlabel metal5 s 15746 5187 16000 6077 6 VSSIO
port 2 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 2 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 2 nsew ground bidirectional
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 2 nsew ground bidirectional
rlabel metal4 s 15746 5167 16000 6097 6 VSSIO
port 2 nsew ground bidirectional
rlabel metal4 s 15746 35157 16000 40000 6 VSSIO
port 2 nsew ground bidirectional
rlabel metal5 s 15746 3977 16000 4867 6 VDDIO
port 3 nsew power bidirectional
rlabel metal5 s 15746 14007 16000 18997 6 VDDIO
port 3 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 3 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 15746 14007 16000 19000 6 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 15746 3957 16000 4887 6 VDDIO
port 3 nsew power bidirectional
rlabel metal5 s 15746 427 16000 1477 6 VCCHIB
port 4 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 4 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 4 nsew power bidirectional
rlabel metal4 s 15746 407 16000 1497 6 VCCHIB
port 4 nsew power bidirectional
rlabel metal5 s 15746 12837 16000 13687 6 VDDIO_Q
port 5 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 5 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 5 nsew power bidirectional
rlabel metal4 s 15746 12817 16000 13707 6 VDDIO_Q
port 5 nsew power bidirectional
rlabel metal5 s 15746 1797 16000 2687 6 VCCD
port 6 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 6 nsew power bidirectional
rlabel metal4 s 15746 1777 16000 2707 6 VCCD
port 6 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 6 nsew power bidirectional
rlabel metal5 s 15746 7368 16000 8017 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 15746 9547 16000 11347 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 11281 16000 11347 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 9547 16000 9613 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 15746 7347 16000 8037 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 15746 10329 16000 10565 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 15746 6397 16000 7047 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 15746 6377 16000 7067 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 15746 11667 16000 12517 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 15746 11647 16000 12537 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 15746 8337 16000 9227 6 VSSD
port 10 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 15746 8317 16000 9247 6 VSSD
port 10 nsew ground bidirectional
rlabel metal5 s 15794 3007 16000 3657 6 VDDA
port 11 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 11 nsew power bidirectional
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 11 nsew power bidirectional
rlabel metal4 s 15794 2987 16000 3677 6 VDDA
port 11 nsew power bidirectional
rlabel metal4 s 0 10625 16000 11221 6 AMUXBUS_A
port 12 nsew signal default
rlabel metal4 s 0 9673 16000 10269 6 AMUXBUS_B
port 13 nsew signal default
<< properties >>
string FIXED_BBOX 0 0 16000 40000
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 192116
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 18226
<< end >>
