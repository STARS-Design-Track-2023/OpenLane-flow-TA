magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1169 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 184 47 214 177
rect 445 47 475 177
rect 529 47 559 177
rect 613 47 643 177
rect 697 47 727 177
rect 805 47 835 177
rect 889 47 919 177
rect 973 47 1003 177
rect 1057 47 1087 177
<< scpmoshvt >>
rect 79 297 109 497
rect 184 297 214 497
rect 372 309 402 497
rect 456 309 486 497
rect 540 309 570 497
rect 624 309 654 497
rect 805 297 835 497
rect 889 297 919 497
rect 973 297 1003 497
rect 1057 297 1087 497
<< ndiff >>
rect 27 106 79 177
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 89 184 177
rect 109 55 119 89
rect 153 55 184 89
rect 109 47 184 55
rect 214 103 266 177
rect 214 69 224 103
rect 258 69 266 103
rect 214 47 266 69
rect 393 129 445 177
rect 393 95 401 129
rect 435 95 445 129
rect 393 47 445 95
rect 475 89 529 177
rect 475 55 485 89
rect 519 55 529 89
rect 475 47 529 55
rect 559 129 613 177
rect 559 95 569 129
rect 603 95 613 129
rect 559 47 613 95
rect 643 89 697 177
rect 643 55 653 89
rect 687 55 697 89
rect 643 47 697 55
rect 727 129 805 177
rect 727 95 749 129
rect 783 95 805 129
rect 727 47 805 95
rect 835 169 889 177
rect 835 135 845 169
rect 879 135 889 169
rect 835 47 889 135
rect 919 89 973 177
rect 919 55 929 89
rect 963 55 973 89
rect 919 47 973 55
rect 1003 169 1057 177
rect 1003 135 1013 169
rect 1047 135 1057 169
rect 1003 47 1057 135
rect 1087 89 1143 177
rect 1087 55 1097 89
rect 1131 55 1143 89
rect 1087 47 1143 55
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 489 184 497
rect 109 455 127 489
rect 161 455 184 489
rect 109 421 184 455
rect 109 387 127 421
rect 161 387 184 421
rect 109 297 184 387
rect 214 477 266 497
rect 214 443 224 477
rect 258 443 266 477
rect 214 409 266 443
rect 214 375 224 409
rect 258 375 266 409
rect 214 297 266 375
rect 320 477 372 497
rect 320 443 328 477
rect 362 443 372 477
rect 320 309 372 443
rect 402 489 456 497
rect 402 455 412 489
rect 446 455 456 489
rect 402 309 456 455
rect 486 477 540 497
rect 486 443 496 477
rect 530 443 540 477
rect 486 309 540 443
rect 570 489 624 497
rect 570 455 580 489
rect 614 455 624 489
rect 570 309 624 455
rect 654 489 805 497
rect 654 387 682 489
rect 784 387 805 489
rect 654 309 805 387
rect 669 297 805 309
rect 835 345 889 497
rect 835 311 845 345
rect 879 311 889 345
rect 835 297 889 311
rect 919 489 973 497
rect 919 455 929 489
rect 963 455 973 489
rect 919 421 973 455
rect 919 387 929 421
rect 963 387 973 421
rect 919 297 973 387
rect 1003 345 1057 497
rect 1003 311 1013 345
rect 1047 311 1057 345
rect 1003 297 1057 311
rect 1087 489 1143 497
rect 1087 455 1097 489
rect 1131 455 1143 489
rect 1087 421 1143 455
rect 1087 387 1097 421
rect 1131 387 1143 421
rect 1087 297 1143 387
<< ndiffc >>
rect 35 72 69 106
rect 119 55 153 89
rect 224 69 258 103
rect 401 95 435 129
rect 485 55 519 89
rect 569 95 603 129
rect 653 55 687 89
rect 749 95 783 129
rect 845 135 879 169
rect 929 55 963 89
rect 1013 135 1047 169
rect 1097 55 1131 89
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 127 455 161 489
rect 127 387 161 421
rect 224 443 258 477
rect 224 375 258 409
rect 328 443 362 477
rect 412 455 446 489
rect 496 443 530 477
rect 580 455 614 489
rect 682 387 784 489
rect 845 311 879 345
rect 929 455 963 489
rect 929 387 963 421
rect 1013 311 1047 345
rect 1097 455 1131 489
rect 1097 387 1131 421
<< poly >>
rect 79 497 109 523
rect 184 497 214 523
rect 372 497 402 523
rect 456 497 486 523
rect 540 497 570 523
rect 624 497 654 523
rect 805 497 835 523
rect 889 497 919 523
rect 973 497 1003 523
rect 1057 497 1087 523
rect 79 265 109 297
rect 184 282 214 297
rect 372 294 402 309
rect 456 294 486 309
rect 540 294 570 309
rect 624 294 654 309
rect 281 282 654 294
rect 79 249 142 265
rect 79 215 98 249
rect 132 215 142 249
rect 79 199 142 215
rect 184 264 654 282
rect 184 252 319 264
rect 805 259 835 297
rect 889 259 919 297
rect 973 259 1003 297
rect 1057 259 1087 297
rect 184 249 260 252
rect 184 215 206 249
rect 240 215 260 249
rect 696 249 762 259
rect 696 222 712 249
rect 184 210 260 215
rect 445 215 712 222
rect 746 215 762 249
rect 184 205 256 210
rect 79 177 109 199
rect 184 177 214 205
rect 445 192 762 215
rect 805 249 1087 259
rect 805 215 833 249
rect 867 215 901 249
rect 935 215 969 249
rect 1003 215 1037 249
rect 1071 215 1087 249
rect 805 205 1087 215
rect 445 177 475 192
rect 529 177 559 192
rect 613 177 643 192
rect 697 177 727 192
rect 805 177 835 205
rect 889 177 919 205
rect 973 177 1003 205
rect 1057 177 1087 205
rect 79 21 109 47
rect 184 21 214 47
rect 445 21 475 47
rect 529 21 559 47
rect 613 21 643 47
rect 697 21 727 47
rect 805 21 835 47
rect 889 21 919 47
rect 973 21 1003 47
rect 1057 21 1087 47
<< polycont >>
rect 98 215 132 249
rect 206 215 240 249
rect 712 215 746 249
rect 833 215 867 249
rect 901 215 935 249
rect 969 215 1003 249
rect 1037 215 1071 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 477 69 493
rect 17 443 35 477
rect 17 409 69 443
rect 17 375 35 409
rect 17 353 69 375
rect 103 489 186 527
rect 103 455 127 489
rect 161 455 186 489
rect 103 421 186 455
rect 103 387 127 421
rect 161 387 186 421
rect 103 369 186 387
rect 220 477 271 493
rect 220 443 224 477
rect 258 443 271 477
rect 220 409 271 443
rect 220 375 224 409
rect 258 375 271 409
rect 313 477 362 493
rect 313 443 328 477
rect 396 489 462 527
rect 396 455 412 489
rect 446 455 462 489
rect 496 477 530 493
rect 313 421 362 443
rect 564 489 630 527
rect 564 455 580 489
rect 614 455 630 489
rect 664 489 1179 493
rect 496 421 530 443
rect 664 421 682 489
rect 313 387 682 421
rect 784 455 929 489
rect 963 455 1097 489
rect 1131 455 1179 489
rect 784 421 1179 455
rect 784 387 929 421
rect 963 387 1097 421
rect 1131 387 1179 421
rect 379 379 1179 387
rect 220 353 271 375
rect 17 255 64 353
rect 17 221 30 255
rect 17 133 64 221
rect 98 249 156 335
rect 220 319 345 353
rect 132 215 156 249
rect 98 153 156 215
rect 190 249 256 285
rect 190 215 206 249
rect 240 215 256 249
rect 190 153 256 215
rect 290 255 345 319
rect 379 311 845 345
rect 879 311 1013 345
rect 1047 311 1179 345
rect 379 289 1179 311
rect 290 249 762 255
rect 290 215 712 249
rect 746 215 762 249
rect 290 205 762 215
rect 796 249 862 255
rect 896 249 1101 255
rect 796 215 833 249
rect 896 221 901 249
rect 867 215 901 221
rect 935 215 969 249
rect 1003 215 1037 249
rect 1071 215 1101 249
rect 796 205 1101 215
rect 17 106 69 133
rect 290 119 345 205
rect 1135 171 1179 289
rect 17 72 35 106
rect 17 56 69 72
rect 103 89 186 119
rect 103 55 119 89
rect 153 55 186 89
rect 103 17 186 55
rect 220 103 345 119
rect 220 69 224 103
rect 258 69 345 103
rect 220 51 345 69
rect 379 131 795 171
rect 379 129 435 131
rect 379 95 401 129
rect 569 129 603 131
rect 379 51 435 95
rect 469 89 535 97
rect 469 55 485 89
rect 519 55 535 89
rect 737 129 795 131
rect 569 55 603 95
rect 637 89 703 97
rect 637 55 653 89
rect 687 55 703 89
rect 469 17 535 55
rect 637 17 703 55
rect 737 95 749 129
rect 783 95 795 129
rect 829 169 1179 171
rect 829 135 845 169
rect 879 135 1013 169
rect 1047 135 1179 169
rect 829 123 1179 135
rect 737 89 795 95
rect 737 55 929 89
rect 963 55 1097 89
rect 1131 55 1147 89
rect 737 51 1147 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 30 221 64 255
rect 862 249 896 255
rect 862 221 867 249
rect 867 221 896 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 17 255 76 261
rect 17 221 30 255
rect 64 252 76 255
rect 850 255 908 261
rect 850 252 862 255
rect 64 224 862 252
rect 64 221 76 224
rect 17 215 76 221
rect 850 221 862 224
rect 896 221 908 255
rect 850 215 908 221
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 122 153 156 187 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 770 289 804 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 678 289 712 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 586 289 620 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 494 289 528 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 402 289 436 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1138 153 1172 187 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1138 221 1172 255 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1138 289 1172 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1046 289 1080 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 954 289 988 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 214 153 248 187 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 122 289 156 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 ebufn_4
rlabel metal1 s 0 -48 1196 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 2956310
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2946864
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
