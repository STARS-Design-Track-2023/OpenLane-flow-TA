magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -66 377 450 897
<< pwell >>
rect -26 -43 410 43
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 384 831
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 831 384 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 384 831
rect 0 791 384 797
rect 0 689 384 763
rect 0 51 384 125
rect 0 17 384 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -23 384 -17
<< labels >>
rlabel metal1 s 0 51 384 125 6 VGND
port 1 nsew ground bidirectional
rlabel metal1 s 0 -23 384 23 8 VNB
port 2 nsew ground bidirectional
rlabel pwell s -26 -43 410 43 8 VNB
port 2 nsew ground bidirectional
rlabel metal1 s 0 791 384 837 6 VPB
port 3 nsew power bidirectional
rlabel nwell s -66 377 450 897 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 0 689 384 763 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 384 814
string LEFclass CORE SPACER
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 91324
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 87792
<< end >>
