magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__nfet_01v8__example_55959141808568  sky130_fd_pr__nfet_01v8__example_55959141808568_0
timestamp 1686671242
transform -1 0 1532 0 1 123
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_0
timestamp 1686671242
transform -1 0 784 0 1 123
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_1
timestamp 1686671242
transform 1 0 840 0 1 123
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_0
timestamp 1686671242
transform 1 0 812 0 1 949
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_1
timestamp 1686671242
transform -1 0 756 0 1 949
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_0
timestamp 1686671242
transform -1 0 4018 0 1 3510
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_1
timestamp 1686671242
transform 1 0 4074 0 1 3510
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808567  sky130_fd_pr__pfet_01v8__example_55959141808567_0
timestamp 1686671242
transform -1 0 4710 0 -1 3710
box -1 0 257 1
<< properties >>
string GDS_END 8176984
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8157906
<< end >>
