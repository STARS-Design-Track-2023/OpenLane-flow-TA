magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< pwell >>
rect 1176 1289 1197 1338
<< locali >>
rect 0 2322 2282 2338
rect 0 2288 80 2322
rect 114 2288 152 2322
rect 186 2288 224 2322
rect 258 2288 296 2322
rect 330 2288 368 2322
rect 402 2288 440 2322
rect 474 2288 512 2322
rect 546 2288 584 2322
rect 618 2288 656 2322
rect 690 2288 728 2322
rect 762 2288 800 2322
rect 834 2288 872 2322
rect 906 2288 944 2322
rect 978 2288 1016 2322
rect 1050 2288 1088 2322
rect 1122 2288 1160 2322
rect 1194 2288 1232 2322
rect 1266 2288 1304 2322
rect 1338 2288 1376 2322
rect 1410 2288 1448 2322
rect 1482 2288 1520 2322
rect 1554 2288 1592 2322
rect 1626 2288 1664 2322
rect 1698 2288 1736 2322
rect 1770 2288 1808 2322
rect 1842 2288 1880 2322
rect 1914 2288 1952 2322
rect 1986 2288 2024 2322
rect 2058 2288 2096 2322
rect 2130 2288 2168 2322
rect 2202 2288 2282 2322
rect 0 2222 2282 2288
rect 0 2188 16 2222
rect 50 2188 2232 2222
rect 2266 2188 2282 2222
rect 0 2150 2282 2188
rect 0 2116 16 2150
rect 50 2116 2232 2150
rect 2266 2116 2282 2150
rect 0 2078 2282 2116
rect 0 2044 16 2078
rect 50 2044 2232 2078
rect 2266 2044 2282 2078
rect 0 2006 2282 2044
rect 0 1972 16 2006
rect 50 1972 2232 2006
rect 2266 1972 2282 2006
rect 0 1934 2282 1972
rect 0 1900 16 1934
rect 50 1900 2232 1934
rect 2266 1900 2282 1934
rect 0 1862 2282 1900
rect 0 1828 16 1862
rect 50 1828 2232 1862
rect 2266 1828 2282 1862
rect 0 1790 2282 1828
rect 0 1756 16 1790
rect 50 1756 2232 1790
rect 2266 1756 2282 1790
rect 0 1718 2282 1756
rect 0 1684 16 1718
rect 50 1684 2232 1718
rect 2266 1684 2282 1718
rect 0 1646 2282 1684
rect 0 1612 16 1646
rect 50 1612 2232 1646
rect 2266 1612 2282 1646
rect 0 1574 2282 1612
rect 0 1540 16 1574
rect 50 1540 2232 1574
rect 2266 1540 2282 1574
rect 0 1502 2282 1540
rect 0 1468 16 1502
rect 50 1468 2232 1502
rect 2266 1468 2282 1502
rect 0 1430 2282 1468
rect 0 1396 16 1430
rect 50 1396 2232 1430
rect 2266 1396 2282 1430
rect 0 1358 2282 1396
rect 0 1324 16 1358
rect 50 1324 2232 1358
rect 2266 1324 2282 1358
rect 0 1286 2282 1324
rect 0 1252 16 1286
rect 50 1252 2232 1286
rect 2266 1252 2282 1286
rect 0 1086 2282 1252
rect 0 1052 16 1086
rect 50 1052 2232 1086
rect 2266 1052 2282 1086
rect 0 1014 2282 1052
rect 0 980 16 1014
rect 50 980 2232 1014
rect 2266 980 2282 1014
rect 0 942 2282 980
rect 0 908 16 942
rect 50 908 2232 942
rect 2266 908 2282 942
rect 0 870 2282 908
rect 0 836 16 870
rect 50 836 2232 870
rect 2266 836 2282 870
rect 0 798 2282 836
rect 0 764 16 798
rect 50 764 2232 798
rect 2266 764 2282 798
rect 0 726 2282 764
rect 0 692 16 726
rect 50 692 2232 726
rect 2266 692 2282 726
rect 0 654 2282 692
rect 0 620 16 654
rect 50 620 2232 654
rect 2266 620 2282 654
rect 0 582 2282 620
rect 0 548 16 582
rect 50 548 2232 582
rect 2266 548 2282 582
rect 0 510 2282 548
rect 0 476 16 510
rect 50 476 2232 510
rect 2266 476 2282 510
rect 0 438 2282 476
rect 0 404 16 438
rect 50 404 2232 438
rect 2266 404 2282 438
rect 0 366 2282 404
rect 0 332 16 366
rect 50 332 2232 366
rect 2266 332 2282 366
rect 0 294 2282 332
rect 0 260 16 294
rect 50 260 2232 294
rect 2266 260 2282 294
rect 0 222 2282 260
rect 0 188 16 222
rect 50 188 2232 222
rect 2266 188 2282 222
rect 0 150 2282 188
rect 0 116 16 150
rect 50 116 2232 150
rect 2266 116 2282 150
rect 0 50 2282 116
rect 0 16 80 50
rect 114 16 152 50
rect 186 16 224 50
rect 258 16 296 50
rect 330 16 368 50
rect 402 16 440 50
rect 474 16 512 50
rect 546 16 584 50
rect 618 16 656 50
rect 690 16 728 50
rect 762 16 800 50
rect 834 16 872 50
rect 906 16 944 50
rect 978 16 1016 50
rect 1050 16 1088 50
rect 1122 16 1160 50
rect 1194 16 1232 50
rect 1266 16 1304 50
rect 1338 16 1376 50
rect 1410 16 1448 50
rect 1482 16 1520 50
rect 1554 16 1592 50
rect 1626 16 1664 50
rect 1698 16 1736 50
rect 1770 16 1808 50
rect 1842 16 1880 50
rect 1914 16 1952 50
rect 1986 16 2024 50
rect 2058 16 2096 50
rect 2130 16 2168 50
rect 2202 16 2282 50
rect 0 0 2282 16
<< viali >>
rect 80 2288 114 2322
rect 152 2288 186 2322
rect 224 2288 258 2322
rect 296 2288 330 2322
rect 368 2288 402 2322
rect 440 2288 474 2322
rect 512 2288 546 2322
rect 584 2288 618 2322
rect 656 2288 690 2322
rect 728 2288 762 2322
rect 800 2288 834 2322
rect 872 2288 906 2322
rect 944 2288 978 2322
rect 1016 2288 1050 2322
rect 1088 2288 1122 2322
rect 1160 2288 1194 2322
rect 1232 2288 1266 2322
rect 1304 2288 1338 2322
rect 1376 2288 1410 2322
rect 1448 2288 1482 2322
rect 1520 2288 1554 2322
rect 1592 2288 1626 2322
rect 1664 2288 1698 2322
rect 1736 2288 1770 2322
rect 1808 2288 1842 2322
rect 1880 2288 1914 2322
rect 1952 2288 1986 2322
rect 2024 2288 2058 2322
rect 2096 2288 2130 2322
rect 2168 2288 2202 2322
rect 16 2188 50 2222
rect 2232 2188 2266 2222
rect 16 2116 50 2150
rect 2232 2116 2266 2150
rect 16 2044 50 2078
rect 2232 2044 2266 2078
rect 16 1972 50 2006
rect 2232 1972 2266 2006
rect 16 1900 50 1934
rect 2232 1900 2266 1934
rect 16 1828 50 1862
rect 2232 1828 2266 1862
rect 16 1756 50 1790
rect 2232 1756 2266 1790
rect 16 1684 50 1718
rect 2232 1684 2266 1718
rect 16 1612 50 1646
rect 2232 1612 2266 1646
rect 16 1540 50 1574
rect 2232 1540 2266 1574
rect 16 1468 50 1502
rect 2232 1468 2266 1502
rect 16 1396 50 1430
rect 2232 1396 2266 1430
rect 16 1324 50 1358
rect 2232 1324 2266 1358
rect 16 1252 50 1286
rect 2232 1252 2266 1286
rect 16 1052 50 1086
rect 2232 1052 2266 1086
rect 16 980 50 1014
rect 2232 980 2266 1014
rect 16 908 50 942
rect 2232 908 2266 942
rect 16 836 50 870
rect 2232 836 2266 870
rect 16 764 50 798
rect 2232 764 2266 798
rect 16 692 50 726
rect 2232 692 2266 726
rect 16 620 50 654
rect 2232 620 2266 654
rect 16 548 50 582
rect 2232 548 2266 582
rect 16 476 50 510
rect 2232 476 2266 510
rect 16 404 50 438
rect 2232 404 2266 438
rect 16 332 50 366
rect 2232 332 2266 366
rect 16 260 50 294
rect 2232 260 2266 294
rect 16 188 50 222
rect 2232 188 2266 222
rect 16 116 50 150
rect 2232 116 2266 150
rect 80 16 114 50
rect 152 16 186 50
rect 224 16 258 50
rect 296 16 330 50
rect 368 16 402 50
rect 440 16 474 50
rect 512 16 546 50
rect 584 16 618 50
rect 656 16 690 50
rect 728 16 762 50
rect 800 16 834 50
rect 872 16 906 50
rect 944 16 978 50
rect 1016 16 1050 50
rect 1088 16 1122 50
rect 1160 16 1194 50
rect 1232 16 1266 50
rect 1304 16 1338 50
rect 1376 16 1410 50
rect 1448 16 1482 50
rect 1520 16 1554 50
rect 1592 16 1626 50
rect 1664 16 1698 50
rect 1736 16 1770 50
rect 1808 16 1842 50
rect 1880 16 1914 50
rect 1952 16 1986 50
rect 2024 16 2058 50
rect 2096 16 2130 50
rect 2168 16 2202 50
<< metal1 >>
rect 0 2331 2282 2338
rect 0 2322 88 2331
rect 0 2288 80 2322
rect 0 2282 88 2288
rect 0 2230 7 2282
rect 59 2279 88 2282
rect 140 2279 152 2331
rect 204 2279 216 2331
rect 268 2279 280 2331
rect 332 2279 344 2331
rect 396 2322 408 2331
rect 460 2322 472 2331
rect 524 2322 536 2331
rect 588 2322 600 2331
rect 652 2322 664 2331
rect 402 2288 408 2322
rect 652 2288 656 2322
rect 396 2279 408 2288
rect 460 2279 472 2288
rect 524 2279 536 2288
rect 588 2279 600 2288
rect 652 2279 664 2288
rect 716 2279 728 2331
rect 780 2279 792 2331
rect 844 2279 856 2331
rect 908 2279 920 2331
rect 972 2322 984 2331
rect 1036 2322 1246 2331
rect 1298 2322 1310 2331
rect 978 2288 984 2322
rect 1050 2288 1088 2322
rect 1122 2288 1160 2322
rect 1194 2288 1232 2322
rect 1298 2288 1304 2322
rect 972 2279 984 2288
rect 1036 2279 1246 2288
rect 1298 2279 1310 2288
rect 1362 2279 1374 2331
rect 1426 2279 1438 2331
rect 1490 2279 1502 2331
rect 1554 2279 1566 2331
rect 1618 2322 1630 2331
rect 1682 2322 1694 2331
rect 1746 2322 1758 2331
rect 1810 2322 1822 2331
rect 1874 2322 1886 2331
rect 1626 2288 1630 2322
rect 1874 2288 1880 2322
rect 1618 2279 1630 2288
rect 1682 2279 1694 2288
rect 1746 2279 1758 2288
rect 1810 2279 1822 2288
rect 1874 2279 1886 2288
rect 1938 2279 1950 2331
rect 2002 2279 2014 2331
rect 2066 2279 2078 2331
rect 2130 2279 2142 2331
rect 2194 2322 2282 2331
rect 2202 2288 2282 2322
rect 2194 2282 2282 2288
rect 2194 2279 2223 2282
rect 59 2272 2223 2279
rect 59 2230 66 2272
rect 0 2222 66 2230
rect 0 2218 16 2222
rect 50 2218 66 2222
rect 0 2166 7 2218
rect 59 2166 66 2218
rect 0 2154 66 2166
rect 0 2102 7 2154
rect 59 2102 66 2154
rect 0 2090 66 2102
rect 0 2038 7 2090
rect 59 2038 66 2090
rect 0 2026 66 2038
rect 0 1974 7 2026
rect 59 1974 66 2026
rect 0 1972 16 1974
rect 50 1972 66 1974
rect 0 1962 66 1972
rect 0 1910 7 1962
rect 59 1910 66 1962
rect 0 1900 16 1910
rect 50 1900 66 1910
rect 0 1898 66 1900
rect 0 1846 7 1898
rect 59 1846 66 1898
rect 0 1834 16 1846
rect 50 1834 66 1846
rect 0 1782 7 1834
rect 59 1782 66 1834
rect 0 1770 16 1782
rect 50 1770 66 1782
rect 0 1718 7 1770
rect 59 1718 66 1770
rect 0 1706 16 1718
rect 50 1706 66 1718
rect 0 1654 7 1706
rect 59 1654 66 1706
rect 0 1646 66 1654
rect 0 1642 16 1646
rect 50 1642 66 1646
rect 0 1590 7 1642
rect 59 1590 66 1642
rect 0 1578 66 1590
rect 0 1526 7 1578
rect 59 1526 66 1578
rect 0 1514 66 1526
rect 0 1462 7 1514
rect 59 1462 66 1514
rect 0 1450 66 1462
rect 0 1398 7 1450
rect 59 1398 66 1450
rect 0 1396 16 1398
rect 50 1396 66 1398
rect 0 1386 66 1396
rect 0 1334 7 1386
rect 59 1334 66 1386
rect 0 1324 16 1334
rect 50 1324 66 1334
rect 0 1322 66 1324
rect 0 1270 7 1322
rect 59 1270 66 1322
rect 0 1252 16 1270
rect 50 1252 66 1270
rect 0 1086 66 1252
rect 0 1068 16 1086
rect 50 1068 66 1086
rect 0 1016 7 1068
rect 59 1016 66 1068
rect 0 1014 66 1016
rect 0 1004 16 1014
rect 50 1004 66 1014
rect 0 952 7 1004
rect 59 952 66 1004
rect 0 942 66 952
rect 0 940 16 942
rect 50 940 66 942
rect 0 888 7 940
rect 59 888 66 940
rect 0 876 66 888
rect 0 824 7 876
rect 59 824 66 876
rect 0 812 66 824
rect 0 760 7 812
rect 59 760 66 812
rect 0 748 66 760
rect 0 696 7 748
rect 59 696 66 748
rect 0 692 16 696
rect 50 692 66 696
rect 0 684 66 692
rect 0 632 7 684
rect 59 632 66 684
rect 0 620 16 632
rect 50 620 66 632
rect 0 568 7 620
rect 59 568 66 620
rect 0 556 16 568
rect 50 556 66 568
rect 0 504 7 556
rect 59 504 66 556
rect 0 492 16 504
rect 50 492 66 504
rect 0 440 7 492
rect 59 440 66 492
rect 0 438 66 440
rect 0 428 16 438
rect 50 428 66 438
rect 0 376 7 428
rect 59 376 66 428
rect 0 366 66 376
rect 0 364 16 366
rect 50 364 66 366
rect 0 312 7 364
rect 59 312 66 364
rect 0 300 66 312
rect 0 248 7 300
rect 59 248 66 300
rect 0 236 66 248
rect 0 184 7 236
rect 59 184 66 236
rect 0 172 66 184
rect 0 120 7 172
rect 59 120 66 172
rect 0 116 16 120
rect 50 116 66 120
rect 0 108 66 116
rect 0 56 7 108
rect 59 66 66 108
rect 100 1201 128 2244
rect 156 1229 184 2272
rect 212 1201 240 2244
rect 268 1229 296 2272
rect 324 1201 352 2244
rect 380 1229 408 2272
rect 436 1201 464 2244
rect 492 1229 520 2272
rect 548 1201 576 2244
rect 604 1229 632 2272
rect 660 1201 688 2244
rect 716 1229 744 2272
rect 772 1201 800 2244
rect 828 1229 856 2272
rect 884 1201 912 2244
rect 940 1229 968 2272
rect 996 1201 1024 2244
rect 1052 1229 1080 2272
rect 1114 2237 1168 2244
rect 1114 2185 1115 2237
rect 1167 2185 1168 2237
rect 1114 2173 1168 2185
rect 1114 2121 1115 2173
rect 1167 2121 1168 2173
rect 1114 2109 1168 2121
rect 1114 2057 1115 2109
rect 1167 2057 1168 2109
rect 1114 2045 1168 2057
rect 1114 1993 1115 2045
rect 1167 1993 1168 2045
rect 1114 1981 1168 1993
rect 1114 1929 1115 1981
rect 1167 1929 1168 1981
rect 1114 1917 1168 1929
rect 1114 1865 1115 1917
rect 1167 1865 1168 1917
rect 1114 1853 1168 1865
rect 1114 1801 1115 1853
rect 1167 1801 1168 1853
rect 1114 1789 1168 1801
rect 1114 1737 1115 1789
rect 1167 1737 1168 1789
rect 1114 1725 1168 1737
rect 1114 1673 1115 1725
rect 1167 1673 1168 1725
rect 1114 1661 1168 1673
rect 1114 1609 1115 1661
rect 1167 1609 1168 1661
rect 1114 1597 1168 1609
rect 1114 1545 1115 1597
rect 1167 1545 1168 1597
rect 1114 1533 1168 1545
rect 1114 1481 1115 1533
rect 1167 1481 1168 1533
rect 1114 1469 1168 1481
rect 1114 1417 1115 1469
rect 1167 1417 1168 1469
rect 1114 1405 1168 1417
rect 1114 1353 1115 1405
rect 1167 1353 1168 1405
rect 1114 1341 1168 1353
rect 1114 1289 1115 1341
rect 1167 1289 1168 1341
rect 1114 1277 1168 1289
rect 1114 1225 1115 1277
rect 1167 1225 1168 1277
rect 1202 1229 1230 2272
rect 1114 1201 1168 1225
rect 1258 1201 1286 2244
rect 1314 1229 1342 2272
rect 1370 1201 1398 2244
rect 1426 1229 1454 2272
rect 1482 1201 1510 2244
rect 1538 1229 1566 2272
rect 1594 1201 1622 2244
rect 1650 1229 1678 2272
rect 1706 1201 1734 2244
rect 1762 1229 1790 2272
rect 1818 1201 1846 2244
rect 1874 1229 1902 2272
rect 1930 1201 1958 2244
rect 1986 1229 2014 2272
rect 2042 1201 2070 2244
rect 2098 1229 2126 2272
rect 2154 1201 2182 2244
rect 100 1195 2182 1201
rect 100 1143 152 1195
rect 204 1143 216 1195
rect 268 1143 280 1195
rect 332 1143 344 1195
rect 396 1143 408 1195
rect 460 1143 472 1195
rect 524 1143 536 1195
rect 588 1143 600 1195
rect 652 1143 664 1195
rect 716 1143 728 1195
rect 780 1143 792 1195
rect 844 1143 856 1195
rect 908 1143 920 1195
rect 972 1143 984 1195
rect 1036 1143 1048 1195
rect 1100 1143 1182 1195
rect 1234 1143 1246 1195
rect 1298 1143 1310 1195
rect 1362 1143 1374 1195
rect 1426 1143 1438 1195
rect 1490 1143 1502 1195
rect 1554 1143 1566 1195
rect 1618 1143 1630 1195
rect 1682 1143 1694 1195
rect 1746 1143 1758 1195
rect 1810 1143 1822 1195
rect 1874 1143 1886 1195
rect 1938 1143 1950 1195
rect 2002 1143 2014 1195
rect 2066 1143 2078 1195
rect 2130 1143 2182 1195
rect 100 1137 2182 1143
rect 100 94 128 1137
rect 156 66 184 1109
rect 212 94 240 1137
rect 268 66 296 1109
rect 324 94 352 1137
rect 380 66 408 1109
rect 436 94 464 1137
rect 492 66 520 1109
rect 548 94 576 1137
rect 604 66 632 1109
rect 660 94 688 1137
rect 716 66 744 1109
rect 772 94 800 1137
rect 828 66 856 1109
rect 884 94 912 1137
rect 940 66 968 1109
rect 996 94 1024 1137
rect 1114 1113 1168 1137
rect 1052 66 1080 1109
rect 1114 1061 1115 1113
rect 1167 1061 1168 1113
rect 1114 1049 1168 1061
rect 1114 997 1115 1049
rect 1167 997 1168 1049
rect 1114 985 1168 997
rect 1114 933 1115 985
rect 1167 933 1168 985
rect 1114 921 1168 933
rect 1114 869 1115 921
rect 1167 869 1168 921
rect 1114 857 1168 869
rect 1114 805 1115 857
rect 1167 805 1168 857
rect 1114 793 1168 805
rect 1114 741 1115 793
rect 1167 741 1168 793
rect 1114 729 1168 741
rect 1114 677 1115 729
rect 1167 677 1168 729
rect 1114 665 1168 677
rect 1114 613 1115 665
rect 1167 613 1168 665
rect 1114 601 1168 613
rect 1114 549 1115 601
rect 1167 549 1168 601
rect 1114 537 1168 549
rect 1114 485 1115 537
rect 1167 485 1168 537
rect 1114 473 1168 485
rect 1114 421 1115 473
rect 1167 421 1168 473
rect 1114 409 1168 421
rect 1114 357 1115 409
rect 1167 357 1168 409
rect 1114 345 1168 357
rect 1114 293 1115 345
rect 1167 293 1168 345
rect 1114 281 1168 293
rect 1114 229 1115 281
rect 1167 229 1168 281
rect 1114 217 1168 229
rect 1114 165 1115 217
rect 1167 165 1168 217
rect 1114 153 1168 165
rect 1114 101 1115 153
rect 1167 101 1168 153
rect 1114 94 1168 101
rect 1202 66 1230 1109
rect 1258 94 1286 1137
rect 1314 66 1342 1109
rect 1370 94 1398 1137
rect 1426 66 1454 1109
rect 1482 94 1510 1137
rect 1538 66 1566 1109
rect 1594 94 1622 1137
rect 1650 66 1678 1109
rect 1706 94 1734 1137
rect 1762 66 1790 1109
rect 1818 94 1846 1137
rect 1874 66 1902 1109
rect 1930 94 1958 1137
rect 1986 66 2014 1109
rect 2042 94 2070 1137
rect 2098 66 2126 1109
rect 2154 94 2182 1137
rect 2216 2230 2223 2272
rect 2275 2230 2282 2282
rect 2216 2222 2282 2230
rect 2216 2218 2232 2222
rect 2266 2218 2282 2222
rect 2216 2166 2223 2218
rect 2275 2166 2282 2218
rect 2216 2154 2282 2166
rect 2216 2102 2223 2154
rect 2275 2102 2282 2154
rect 2216 2090 2282 2102
rect 2216 2038 2223 2090
rect 2275 2038 2282 2090
rect 2216 2026 2282 2038
rect 2216 1974 2223 2026
rect 2275 1974 2282 2026
rect 2216 1972 2232 1974
rect 2266 1972 2282 1974
rect 2216 1962 2282 1972
rect 2216 1910 2223 1962
rect 2275 1910 2282 1962
rect 2216 1900 2232 1910
rect 2266 1900 2282 1910
rect 2216 1898 2282 1900
rect 2216 1846 2223 1898
rect 2275 1846 2282 1898
rect 2216 1834 2232 1846
rect 2266 1834 2282 1846
rect 2216 1782 2223 1834
rect 2275 1782 2282 1834
rect 2216 1770 2232 1782
rect 2266 1770 2282 1782
rect 2216 1718 2223 1770
rect 2275 1718 2282 1770
rect 2216 1706 2232 1718
rect 2266 1706 2282 1718
rect 2216 1654 2223 1706
rect 2275 1654 2282 1706
rect 2216 1646 2282 1654
rect 2216 1642 2232 1646
rect 2266 1642 2282 1646
rect 2216 1590 2223 1642
rect 2275 1590 2282 1642
rect 2216 1578 2282 1590
rect 2216 1526 2223 1578
rect 2275 1526 2282 1578
rect 2216 1514 2282 1526
rect 2216 1462 2223 1514
rect 2275 1462 2282 1514
rect 2216 1450 2282 1462
rect 2216 1398 2223 1450
rect 2275 1398 2282 1450
rect 2216 1396 2232 1398
rect 2266 1396 2282 1398
rect 2216 1386 2282 1396
rect 2216 1334 2223 1386
rect 2275 1334 2282 1386
rect 2216 1324 2232 1334
rect 2266 1324 2282 1334
rect 2216 1322 2282 1324
rect 2216 1270 2223 1322
rect 2275 1270 2282 1322
rect 2216 1252 2232 1270
rect 2266 1252 2282 1270
rect 2216 1086 2282 1252
rect 2216 1068 2232 1086
rect 2266 1068 2282 1086
rect 2216 1016 2223 1068
rect 2275 1016 2282 1068
rect 2216 1014 2282 1016
rect 2216 1004 2232 1014
rect 2266 1004 2282 1014
rect 2216 952 2223 1004
rect 2275 952 2282 1004
rect 2216 942 2282 952
rect 2216 940 2232 942
rect 2266 940 2282 942
rect 2216 888 2223 940
rect 2275 888 2282 940
rect 2216 876 2282 888
rect 2216 824 2223 876
rect 2275 824 2282 876
rect 2216 812 2282 824
rect 2216 760 2223 812
rect 2275 760 2282 812
rect 2216 748 2282 760
rect 2216 696 2223 748
rect 2275 696 2282 748
rect 2216 692 2232 696
rect 2266 692 2282 696
rect 2216 684 2282 692
rect 2216 632 2223 684
rect 2275 632 2282 684
rect 2216 620 2232 632
rect 2266 620 2282 632
rect 2216 568 2223 620
rect 2275 568 2282 620
rect 2216 556 2232 568
rect 2266 556 2282 568
rect 2216 504 2223 556
rect 2275 504 2282 556
rect 2216 492 2232 504
rect 2266 492 2282 504
rect 2216 440 2223 492
rect 2275 440 2282 492
rect 2216 438 2282 440
rect 2216 428 2232 438
rect 2266 428 2282 438
rect 2216 376 2223 428
rect 2275 376 2282 428
rect 2216 366 2282 376
rect 2216 364 2232 366
rect 2266 364 2282 366
rect 2216 312 2223 364
rect 2275 312 2282 364
rect 2216 300 2282 312
rect 2216 248 2223 300
rect 2275 248 2282 300
rect 2216 236 2282 248
rect 2216 184 2223 236
rect 2275 184 2282 236
rect 2216 172 2282 184
rect 2216 120 2223 172
rect 2275 120 2282 172
rect 2216 116 2232 120
rect 2266 116 2282 120
rect 2216 108 2282 116
rect 2216 66 2223 108
rect 59 59 2223 66
rect 59 56 88 59
rect 0 50 88 56
rect 0 16 80 50
rect 0 7 88 16
rect 140 7 152 59
rect 204 7 216 59
rect 268 7 280 59
rect 332 7 344 59
rect 396 50 408 59
rect 460 50 472 59
rect 524 50 536 59
rect 588 50 600 59
rect 652 50 664 59
rect 402 16 408 50
rect 652 16 656 50
rect 396 7 408 16
rect 460 7 472 16
rect 524 7 536 16
rect 588 7 600 16
rect 652 7 664 16
rect 716 7 728 59
rect 780 7 792 59
rect 844 7 856 59
rect 908 7 920 59
rect 972 50 984 59
rect 1036 50 1246 59
rect 1298 50 1310 59
rect 978 16 984 50
rect 1050 16 1088 50
rect 1122 16 1160 50
rect 1194 16 1232 50
rect 1298 16 1304 50
rect 972 7 984 16
rect 1036 7 1246 16
rect 1298 7 1310 16
rect 1362 7 1374 59
rect 1426 7 1438 59
rect 1490 7 1502 59
rect 1554 7 1566 59
rect 1618 50 1630 59
rect 1682 50 1694 59
rect 1746 50 1758 59
rect 1810 50 1822 59
rect 1874 50 1886 59
rect 1626 16 1630 50
rect 1874 16 1880 50
rect 1618 7 1630 16
rect 1682 7 1694 16
rect 1746 7 1758 16
rect 1810 7 1822 16
rect 1874 7 1886 16
rect 1938 7 1950 59
rect 2002 7 2014 59
rect 2066 7 2078 59
rect 2130 7 2142 59
rect 2194 56 2223 59
rect 2275 56 2282 108
rect 2194 50 2282 56
rect 2202 16 2282 50
rect 2194 7 2282 16
rect 0 0 2282 7
<< via1 >>
rect 88 2322 140 2331
rect 88 2288 114 2322
rect 114 2288 140 2322
rect 7 2230 59 2282
rect 88 2279 140 2288
rect 152 2322 204 2331
rect 152 2288 186 2322
rect 186 2288 204 2322
rect 152 2279 204 2288
rect 216 2322 268 2331
rect 216 2288 224 2322
rect 224 2288 258 2322
rect 258 2288 268 2322
rect 216 2279 268 2288
rect 280 2322 332 2331
rect 280 2288 296 2322
rect 296 2288 330 2322
rect 330 2288 332 2322
rect 280 2279 332 2288
rect 344 2322 396 2331
rect 408 2322 460 2331
rect 472 2322 524 2331
rect 536 2322 588 2331
rect 600 2322 652 2331
rect 664 2322 716 2331
rect 344 2288 368 2322
rect 368 2288 396 2322
rect 408 2288 440 2322
rect 440 2288 460 2322
rect 472 2288 474 2322
rect 474 2288 512 2322
rect 512 2288 524 2322
rect 536 2288 546 2322
rect 546 2288 584 2322
rect 584 2288 588 2322
rect 600 2288 618 2322
rect 618 2288 652 2322
rect 664 2288 690 2322
rect 690 2288 716 2322
rect 344 2279 396 2288
rect 408 2279 460 2288
rect 472 2279 524 2288
rect 536 2279 588 2288
rect 600 2279 652 2288
rect 664 2279 716 2288
rect 728 2322 780 2331
rect 728 2288 762 2322
rect 762 2288 780 2322
rect 728 2279 780 2288
rect 792 2322 844 2331
rect 792 2288 800 2322
rect 800 2288 834 2322
rect 834 2288 844 2322
rect 792 2279 844 2288
rect 856 2322 908 2331
rect 856 2288 872 2322
rect 872 2288 906 2322
rect 906 2288 908 2322
rect 856 2279 908 2288
rect 920 2322 972 2331
rect 984 2322 1036 2331
rect 1246 2322 1298 2331
rect 1310 2322 1362 2331
rect 920 2288 944 2322
rect 944 2288 972 2322
rect 984 2288 1016 2322
rect 1016 2288 1036 2322
rect 1246 2288 1266 2322
rect 1266 2288 1298 2322
rect 1310 2288 1338 2322
rect 1338 2288 1362 2322
rect 920 2279 972 2288
rect 984 2279 1036 2288
rect 1246 2279 1298 2288
rect 1310 2279 1362 2288
rect 1374 2322 1426 2331
rect 1374 2288 1376 2322
rect 1376 2288 1410 2322
rect 1410 2288 1426 2322
rect 1374 2279 1426 2288
rect 1438 2322 1490 2331
rect 1438 2288 1448 2322
rect 1448 2288 1482 2322
rect 1482 2288 1490 2322
rect 1438 2279 1490 2288
rect 1502 2322 1554 2331
rect 1502 2288 1520 2322
rect 1520 2288 1554 2322
rect 1502 2279 1554 2288
rect 1566 2322 1618 2331
rect 1630 2322 1682 2331
rect 1694 2322 1746 2331
rect 1758 2322 1810 2331
rect 1822 2322 1874 2331
rect 1886 2322 1938 2331
rect 1566 2288 1592 2322
rect 1592 2288 1618 2322
rect 1630 2288 1664 2322
rect 1664 2288 1682 2322
rect 1694 2288 1698 2322
rect 1698 2288 1736 2322
rect 1736 2288 1746 2322
rect 1758 2288 1770 2322
rect 1770 2288 1808 2322
rect 1808 2288 1810 2322
rect 1822 2288 1842 2322
rect 1842 2288 1874 2322
rect 1886 2288 1914 2322
rect 1914 2288 1938 2322
rect 1566 2279 1618 2288
rect 1630 2279 1682 2288
rect 1694 2279 1746 2288
rect 1758 2279 1810 2288
rect 1822 2279 1874 2288
rect 1886 2279 1938 2288
rect 1950 2322 2002 2331
rect 1950 2288 1952 2322
rect 1952 2288 1986 2322
rect 1986 2288 2002 2322
rect 1950 2279 2002 2288
rect 2014 2322 2066 2331
rect 2014 2288 2024 2322
rect 2024 2288 2058 2322
rect 2058 2288 2066 2322
rect 2014 2279 2066 2288
rect 2078 2322 2130 2331
rect 2078 2288 2096 2322
rect 2096 2288 2130 2322
rect 2078 2279 2130 2288
rect 2142 2322 2194 2331
rect 2142 2288 2168 2322
rect 2168 2288 2194 2322
rect 2142 2279 2194 2288
rect 7 2188 16 2218
rect 16 2188 50 2218
rect 50 2188 59 2218
rect 7 2166 59 2188
rect 7 2150 59 2154
rect 7 2116 16 2150
rect 16 2116 50 2150
rect 50 2116 59 2150
rect 7 2102 59 2116
rect 7 2078 59 2090
rect 7 2044 16 2078
rect 16 2044 50 2078
rect 50 2044 59 2078
rect 7 2038 59 2044
rect 7 2006 59 2026
rect 7 1974 16 2006
rect 16 1974 50 2006
rect 50 1974 59 2006
rect 7 1934 59 1962
rect 7 1910 16 1934
rect 16 1910 50 1934
rect 50 1910 59 1934
rect 7 1862 59 1898
rect 7 1846 16 1862
rect 16 1846 50 1862
rect 50 1846 59 1862
rect 7 1828 16 1834
rect 16 1828 50 1834
rect 50 1828 59 1834
rect 7 1790 59 1828
rect 7 1782 16 1790
rect 16 1782 50 1790
rect 50 1782 59 1790
rect 7 1756 16 1770
rect 16 1756 50 1770
rect 50 1756 59 1770
rect 7 1718 59 1756
rect 7 1684 16 1706
rect 16 1684 50 1706
rect 50 1684 59 1706
rect 7 1654 59 1684
rect 7 1612 16 1642
rect 16 1612 50 1642
rect 50 1612 59 1642
rect 7 1590 59 1612
rect 7 1574 59 1578
rect 7 1540 16 1574
rect 16 1540 50 1574
rect 50 1540 59 1574
rect 7 1526 59 1540
rect 7 1502 59 1514
rect 7 1468 16 1502
rect 16 1468 50 1502
rect 50 1468 59 1502
rect 7 1462 59 1468
rect 7 1430 59 1450
rect 7 1398 16 1430
rect 16 1398 50 1430
rect 50 1398 59 1430
rect 7 1358 59 1386
rect 7 1334 16 1358
rect 16 1334 50 1358
rect 50 1334 59 1358
rect 7 1286 59 1322
rect 7 1270 16 1286
rect 16 1270 50 1286
rect 50 1270 59 1286
rect 7 1052 16 1068
rect 16 1052 50 1068
rect 50 1052 59 1068
rect 7 1016 59 1052
rect 7 980 16 1004
rect 16 980 50 1004
rect 50 980 59 1004
rect 7 952 59 980
rect 7 908 16 940
rect 16 908 50 940
rect 50 908 59 940
rect 7 888 59 908
rect 7 870 59 876
rect 7 836 16 870
rect 16 836 50 870
rect 50 836 59 870
rect 7 824 59 836
rect 7 798 59 812
rect 7 764 16 798
rect 16 764 50 798
rect 50 764 59 798
rect 7 760 59 764
rect 7 726 59 748
rect 7 696 16 726
rect 16 696 50 726
rect 50 696 59 726
rect 7 654 59 684
rect 7 632 16 654
rect 16 632 50 654
rect 50 632 59 654
rect 7 582 59 620
rect 7 568 16 582
rect 16 568 50 582
rect 50 568 59 582
rect 7 548 16 556
rect 16 548 50 556
rect 50 548 59 556
rect 7 510 59 548
rect 7 504 16 510
rect 16 504 50 510
rect 50 504 59 510
rect 7 476 16 492
rect 16 476 50 492
rect 50 476 59 492
rect 7 440 59 476
rect 7 404 16 428
rect 16 404 50 428
rect 50 404 59 428
rect 7 376 59 404
rect 7 332 16 364
rect 16 332 50 364
rect 50 332 59 364
rect 7 312 59 332
rect 7 294 59 300
rect 7 260 16 294
rect 16 260 50 294
rect 50 260 59 294
rect 7 248 59 260
rect 7 222 59 236
rect 7 188 16 222
rect 16 188 50 222
rect 50 188 59 222
rect 7 184 59 188
rect 7 150 59 172
rect 7 120 16 150
rect 16 120 50 150
rect 50 120 59 150
rect 7 56 59 108
rect 1115 2185 1167 2237
rect 1115 2121 1167 2173
rect 1115 2057 1167 2109
rect 1115 1993 1167 2045
rect 1115 1929 1167 1981
rect 1115 1865 1167 1917
rect 1115 1801 1167 1853
rect 1115 1737 1167 1789
rect 1115 1673 1167 1725
rect 1115 1609 1167 1661
rect 1115 1545 1167 1597
rect 1115 1481 1167 1533
rect 1115 1417 1167 1469
rect 1115 1353 1167 1405
rect 1115 1289 1167 1341
rect 1115 1225 1167 1277
rect 152 1143 204 1195
rect 216 1143 268 1195
rect 280 1143 332 1195
rect 344 1143 396 1195
rect 408 1143 460 1195
rect 472 1143 524 1195
rect 536 1143 588 1195
rect 600 1143 652 1195
rect 664 1143 716 1195
rect 728 1143 780 1195
rect 792 1143 844 1195
rect 856 1143 908 1195
rect 920 1143 972 1195
rect 984 1143 1036 1195
rect 1048 1143 1100 1195
rect 1182 1143 1234 1195
rect 1246 1143 1298 1195
rect 1310 1143 1362 1195
rect 1374 1143 1426 1195
rect 1438 1143 1490 1195
rect 1502 1143 1554 1195
rect 1566 1143 1618 1195
rect 1630 1143 1682 1195
rect 1694 1143 1746 1195
rect 1758 1143 1810 1195
rect 1822 1143 1874 1195
rect 1886 1143 1938 1195
rect 1950 1143 2002 1195
rect 2014 1143 2066 1195
rect 2078 1143 2130 1195
rect 1115 1061 1167 1113
rect 1115 997 1167 1049
rect 1115 933 1167 985
rect 1115 869 1167 921
rect 1115 805 1167 857
rect 1115 741 1167 793
rect 1115 677 1167 729
rect 1115 613 1167 665
rect 1115 549 1167 601
rect 1115 485 1167 537
rect 1115 421 1167 473
rect 1115 357 1167 409
rect 1115 293 1167 345
rect 1115 229 1167 281
rect 1115 165 1167 217
rect 1115 101 1167 153
rect 2223 2230 2275 2282
rect 2223 2188 2232 2218
rect 2232 2188 2266 2218
rect 2266 2188 2275 2218
rect 2223 2166 2275 2188
rect 2223 2150 2275 2154
rect 2223 2116 2232 2150
rect 2232 2116 2266 2150
rect 2266 2116 2275 2150
rect 2223 2102 2275 2116
rect 2223 2078 2275 2090
rect 2223 2044 2232 2078
rect 2232 2044 2266 2078
rect 2266 2044 2275 2078
rect 2223 2038 2275 2044
rect 2223 2006 2275 2026
rect 2223 1974 2232 2006
rect 2232 1974 2266 2006
rect 2266 1974 2275 2006
rect 2223 1934 2275 1962
rect 2223 1910 2232 1934
rect 2232 1910 2266 1934
rect 2266 1910 2275 1934
rect 2223 1862 2275 1898
rect 2223 1846 2232 1862
rect 2232 1846 2266 1862
rect 2266 1846 2275 1862
rect 2223 1828 2232 1834
rect 2232 1828 2266 1834
rect 2266 1828 2275 1834
rect 2223 1790 2275 1828
rect 2223 1782 2232 1790
rect 2232 1782 2266 1790
rect 2266 1782 2275 1790
rect 2223 1756 2232 1770
rect 2232 1756 2266 1770
rect 2266 1756 2275 1770
rect 2223 1718 2275 1756
rect 2223 1684 2232 1706
rect 2232 1684 2266 1706
rect 2266 1684 2275 1706
rect 2223 1654 2275 1684
rect 2223 1612 2232 1642
rect 2232 1612 2266 1642
rect 2266 1612 2275 1642
rect 2223 1590 2275 1612
rect 2223 1574 2275 1578
rect 2223 1540 2232 1574
rect 2232 1540 2266 1574
rect 2266 1540 2275 1574
rect 2223 1526 2275 1540
rect 2223 1502 2275 1514
rect 2223 1468 2232 1502
rect 2232 1468 2266 1502
rect 2266 1468 2275 1502
rect 2223 1462 2275 1468
rect 2223 1430 2275 1450
rect 2223 1398 2232 1430
rect 2232 1398 2266 1430
rect 2266 1398 2275 1430
rect 2223 1358 2275 1386
rect 2223 1334 2232 1358
rect 2232 1334 2266 1358
rect 2266 1334 2275 1358
rect 2223 1286 2275 1322
rect 2223 1270 2232 1286
rect 2232 1270 2266 1286
rect 2266 1270 2275 1286
rect 2223 1052 2232 1068
rect 2232 1052 2266 1068
rect 2266 1052 2275 1068
rect 2223 1016 2275 1052
rect 2223 980 2232 1004
rect 2232 980 2266 1004
rect 2266 980 2275 1004
rect 2223 952 2275 980
rect 2223 908 2232 940
rect 2232 908 2266 940
rect 2266 908 2275 940
rect 2223 888 2275 908
rect 2223 870 2275 876
rect 2223 836 2232 870
rect 2232 836 2266 870
rect 2266 836 2275 870
rect 2223 824 2275 836
rect 2223 798 2275 812
rect 2223 764 2232 798
rect 2232 764 2266 798
rect 2266 764 2275 798
rect 2223 760 2275 764
rect 2223 726 2275 748
rect 2223 696 2232 726
rect 2232 696 2266 726
rect 2266 696 2275 726
rect 2223 654 2275 684
rect 2223 632 2232 654
rect 2232 632 2266 654
rect 2266 632 2275 654
rect 2223 582 2275 620
rect 2223 568 2232 582
rect 2232 568 2266 582
rect 2266 568 2275 582
rect 2223 548 2232 556
rect 2232 548 2266 556
rect 2266 548 2275 556
rect 2223 510 2275 548
rect 2223 504 2232 510
rect 2232 504 2266 510
rect 2266 504 2275 510
rect 2223 476 2232 492
rect 2232 476 2266 492
rect 2266 476 2275 492
rect 2223 440 2275 476
rect 2223 404 2232 428
rect 2232 404 2266 428
rect 2266 404 2275 428
rect 2223 376 2275 404
rect 2223 332 2232 364
rect 2232 332 2266 364
rect 2266 332 2275 364
rect 2223 312 2275 332
rect 2223 294 2275 300
rect 2223 260 2232 294
rect 2232 260 2266 294
rect 2266 260 2275 294
rect 2223 248 2275 260
rect 2223 222 2275 236
rect 2223 188 2232 222
rect 2232 188 2266 222
rect 2266 188 2275 222
rect 2223 184 2275 188
rect 2223 150 2275 172
rect 2223 120 2232 150
rect 2232 120 2266 150
rect 2266 120 2275 150
rect 88 50 140 59
rect 88 16 114 50
rect 114 16 140 50
rect 88 7 140 16
rect 152 50 204 59
rect 152 16 186 50
rect 186 16 204 50
rect 152 7 204 16
rect 216 50 268 59
rect 216 16 224 50
rect 224 16 258 50
rect 258 16 268 50
rect 216 7 268 16
rect 280 50 332 59
rect 280 16 296 50
rect 296 16 330 50
rect 330 16 332 50
rect 280 7 332 16
rect 344 50 396 59
rect 408 50 460 59
rect 472 50 524 59
rect 536 50 588 59
rect 600 50 652 59
rect 664 50 716 59
rect 344 16 368 50
rect 368 16 396 50
rect 408 16 440 50
rect 440 16 460 50
rect 472 16 474 50
rect 474 16 512 50
rect 512 16 524 50
rect 536 16 546 50
rect 546 16 584 50
rect 584 16 588 50
rect 600 16 618 50
rect 618 16 652 50
rect 664 16 690 50
rect 690 16 716 50
rect 344 7 396 16
rect 408 7 460 16
rect 472 7 524 16
rect 536 7 588 16
rect 600 7 652 16
rect 664 7 716 16
rect 728 50 780 59
rect 728 16 762 50
rect 762 16 780 50
rect 728 7 780 16
rect 792 50 844 59
rect 792 16 800 50
rect 800 16 834 50
rect 834 16 844 50
rect 792 7 844 16
rect 856 50 908 59
rect 856 16 872 50
rect 872 16 906 50
rect 906 16 908 50
rect 856 7 908 16
rect 920 50 972 59
rect 984 50 1036 59
rect 1246 50 1298 59
rect 1310 50 1362 59
rect 920 16 944 50
rect 944 16 972 50
rect 984 16 1016 50
rect 1016 16 1036 50
rect 1246 16 1266 50
rect 1266 16 1298 50
rect 1310 16 1338 50
rect 1338 16 1362 50
rect 920 7 972 16
rect 984 7 1036 16
rect 1246 7 1298 16
rect 1310 7 1362 16
rect 1374 50 1426 59
rect 1374 16 1376 50
rect 1376 16 1410 50
rect 1410 16 1426 50
rect 1374 7 1426 16
rect 1438 50 1490 59
rect 1438 16 1448 50
rect 1448 16 1482 50
rect 1482 16 1490 50
rect 1438 7 1490 16
rect 1502 50 1554 59
rect 1502 16 1520 50
rect 1520 16 1554 50
rect 1502 7 1554 16
rect 1566 50 1618 59
rect 1630 50 1682 59
rect 1694 50 1746 59
rect 1758 50 1810 59
rect 1822 50 1874 59
rect 1886 50 1938 59
rect 1566 16 1592 50
rect 1592 16 1618 50
rect 1630 16 1664 50
rect 1664 16 1682 50
rect 1694 16 1698 50
rect 1698 16 1736 50
rect 1736 16 1746 50
rect 1758 16 1770 50
rect 1770 16 1808 50
rect 1808 16 1810 50
rect 1822 16 1842 50
rect 1842 16 1874 50
rect 1886 16 1914 50
rect 1914 16 1938 50
rect 1566 7 1618 16
rect 1630 7 1682 16
rect 1694 7 1746 16
rect 1758 7 1810 16
rect 1822 7 1874 16
rect 1886 7 1938 16
rect 1950 50 2002 59
rect 1950 16 1952 50
rect 1952 16 1986 50
rect 1986 16 2002 50
rect 1950 7 2002 16
rect 2014 50 2066 59
rect 2014 16 2024 50
rect 2024 16 2058 50
rect 2058 16 2066 50
rect 2014 7 2066 16
rect 2078 50 2130 59
rect 2078 16 2096 50
rect 2096 16 2130 50
rect 2078 7 2130 16
rect 2142 50 2194 59
rect 2223 56 2275 108
rect 2142 16 2168 50
rect 2168 16 2194 50
rect 2142 7 2194 16
<< metal2 >>
rect 0 2331 1086 2338
rect 0 2282 88 2331
rect 0 2230 7 2282
rect 59 2279 88 2282
rect 140 2279 152 2331
rect 204 2279 216 2331
rect 268 2279 280 2331
rect 332 2279 344 2331
rect 396 2279 408 2331
rect 460 2279 472 2331
rect 524 2279 536 2331
rect 588 2279 600 2331
rect 652 2279 664 2331
rect 716 2279 728 2331
rect 780 2279 792 2331
rect 844 2279 856 2331
rect 908 2279 920 2331
rect 972 2279 984 2331
rect 1036 2279 1086 2331
rect 59 2272 1086 2279
rect 59 2230 66 2272
rect 1114 2244 1168 2338
rect 1196 2331 2282 2338
rect 1196 2279 1246 2331
rect 1298 2279 1310 2331
rect 1362 2279 1374 2331
rect 1426 2279 1438 2331
rect 1490 2279 1502 2331
rect 1554 2279 1566 2331
rect 1618 2279 1630 2331
rect 1682 2279 1694 2331
rect 1746 2279 1758 2331
rect 1810 2279 1822 2331
rect 1874 2279 1886 2331
rect 1938 2279 1950 2331
rect 2002 2279 2014 2331
rect 2066 2279 2078 2331
rect 2130 2279 2142 2331
rect 2194 2282 2282 2331
rect 2194 2279 2223 2282
rect 1196 2272 2223 2279
rect 0 2218 66 2230
rect 0 2166 7 2218
rect 59 2188 66 2218
rect 94 2237 2188 2244
rect 94 2216 1115 2237
rect 59 2166 1086 2188
rect 0 2160 1086 2166
rect 1114 2185 1115 2216
rect 1167 2216 2188 2237
rect 2216 2230 2223 2272
rect 2275 2230 2282 2282
rect 2216 2218 2282 2230
rect 1167 2185 1168 2216
rect 2216 2188 2223 2218
rect 1114 2173 1168 2185
rect 0 2154 66 2160
rect 0 2102 7 2154
rect 59 2102 66 2154
rect 1114 2132 1115 2173
rect 94 2121 1115 2132
rect 1167 2132 1168 2173
rect 1196 2166 2223 2188
rect 2275 2166 2282 2218
rect 1196 2160 2282 2166
rect 2216 2154 2282 2160
rect 1167 2121 2188 2132
rect 94 2109 2188 2121
rect 94 2104 1115 2109
rect 0 2090 66 2102
rect 0 2038 7 2090
rect 59 2076 66 2090
rect 59 2048 1086 2076
rect 1114 2057 1115 2104
rect 1167 2104 2188 2109
rect 1167 2057 1168 2104
rect 2216 2102 2223 2154
rect 2275 2102 2282 2154
rect 2216 2090 2282 2102
rect 2216 2076 2223 2090
rect 59 2038 66 2048
rect 0 2026 66 2038
rect 0 1974 7 2026
rect 59 1974 66 2026
rect 1114 2045 1168 2057
rect 1196 2048 2223 2076
rect 1114 2020 1115 2045
rect 94 1993 1115 2020
rect 1167 2020 1168 2045
rect 2216 2038 2223 2048
rect 2275 2038 2282 2090
rect 2216 2026 2282 2038
rect 1167 1993 2188 2020
rect 94 1992 2188 1993
rect 0 1964 66 1974
rect 1114 1981 1168 1992
rect 0 1962 1086 1964
rect 0 1910 7 1962
rect 59 1936 1086 1962
rect 59 1910 66 1936
rect 0 1898 66 1910
rect 1114 1929 1115 1981
rect 1167 1929 1168 1981
rect 2216 1974 2223 2026
rect 2275 1974 2282 2026
rect 2216 1964 2282 1974
rect 1196 1962 2282 1964
rect 1196 1936 2223 1962
rect 1114 1917 1168 1929
rect 1114 1908 1115 1917
rect 0 1846 7 1898
rect 59 1852 66 1898
rect 94 1880 1115 1908
rect 1114 1865 1115 1880
rect 1167 1908 1168 1917
rect 2216 1910 2223 1936
rect 2275 1910 2282 1962
rect 1167 1880 2188 1908
rect 2216 1898 2282 1910
rect 1167 1865 1168 1880
rect 1114 1853 1168 1865
rect 59 1846 1086 1852
rect 0 1834 1086 1846
rect 0 1782 7 1834
rect 59 1824 1086 1834
rect 59 1782 66 1824
rect 1114 1801 1115 1853
rect 1167 1801 1168 1853
rect 2216 1852 2223 1898
rect 1196 1846 2223 1852
rect 2275 1846 2282 1898
rect 1196 1834 2282 1846
rect 1196 1824 2223 1834
rect 1114 1796 1168 1801
rect 0 1770 66 1782
rect 0 1718 7 1770
rect 59 1740 66 1770
rect 94 1789 2188 1796
rect 94 1768 1115 1789
rect 59 1718 1086 1740
rect 0 1712 1086 1718
rect 1114 1737 1115 1768
rect 1167 1768 2188 1789
rect 2216 1782 2223 1824
rect 2275 1782 2282 1834
rect 2216 1770 2282 1782
rect 1167 1737 1168 1768
rect 2216 1740 2223 1770
rect 1114 1725 1168 1737
rect 0 1706 66 1712
rect 0 1654 7 1706
rect 59 1654 66 1706
rect 1114 1684 1115 1725
rect 94 1673 1115 1684
rect 1167 1684 1168 1725
rect 1196 1718 2223 1740
rect 2275 1718 2282 1770
rect 1196 1712 2282 1718
rect 2216 1706 2282 1712
rect 1167 1673 2188 1684
rect 94 1661 2188 1673
rect 94 1656 1115 1661
rect 0 1642 66 1654
rect 0 1590 7 1642
rect 59 1628 66 1642
rect 59 1600 1086 1628
rect 1114 1609 1115 1656
rect 1167 1656 2188 1661
rect 1167 1609 1168 1656
rect 2216 1654 2223 1706
rect 2275 1654 2282 1706
rect 2216 1642 2282 1654
rect 2216 1628 2223 1642
rect 59 1590 66 1600
rect 0 1578 66 1590
rect 0 1526 7 1578
rect 59 1526 66 1578
rect 1114 1597 1168 1609
rect 1196 1600 2223 1628
rect 1114 1572 1115 1597
rect 94 1545 1115 1572
rect 1167 1572 1168 1597
rect 2216 1590 2223 1600
rect 2275 1590 2282 1642
rect 2216 1578 2282 1590
rect 1167 1545 2188 1572
rect 94 1544 2188 1545
rect 0 1516 66 1526
rect 1114 1533 1168 1544
rect 0 1514 1086 1516
rect 0 1462 7 1514
rect 59 1488 1086 1514
rect 59 1462 66 1488
rect 0 1450 66 1462
rect 1114 1481 1115 1533
rect 1167 1481 1168 1533
rect 2216 1526 2223 1578
rect 2275 1526 2282 1578
rect 2216 1516 2282 1526
rect 1196 1514 2282 1516
rect 1196 1488 2223 1514
rect 1114 1469 1168 1481
rect 1114 1460 1115 1469
rect 0 1398 7 1450
rect 59 1404 66 1450
rect 94 1432 1115 1460
rect 1114 1417 1115 1432
rect 1167 1460 1168 1469
rect 2216 1462 2223 1488
rect 2275 1462 2282 1514
rect 1167 1432 2188 1460
rect 2216 1450 2282 1462
rect 1167 1417 1168 1432
rect 1114 1405 1168 1417
rect 59 1398 1086 1404
rect 0 1386 1086 1398
rect 0 1334 7 1386
rect 59 1376 1086 1386
rect 59 1334 66 1376
rect 1114 1353 1115 1405
rect 1167 1353 1168 1405
rect 2216 1404 2223 1450
rect 1196 1398 2223 1404
rect 2275 1398 2282 1450
rect 1196 1386 2282 1398
rect 1196 1376 2223 1386
rect 1114 1348 1168 1353
rect 0 1322 66 1334
rect 0 1270 7 1322
rect 59 1292 66 1322
rect 94 1341 2188 1348
rect 94 1320 1115 1341
rect 59 1270 1086 1292
rect 0 1224 1086 1270
rect 1114 1289 1115 1320
rect 1167 1320 2188 1341
rect 2216 1334 2223 1376
rect 2275 1334 2282 1386
rect 2216 1322 2282 1334
rect 1167 1289 1168 1320
rect 2216 1292 2223 1322
rect 1114 1277 1168 1289
rect 1114 1225 1115 1277
rect 1167 1225 1168 1277
rect 1114 1196 1168 1225
rect 1196 1270 2223 1292
rect 2275 1270 2282 1322
rect 1196 1224 2282 1270
rect 0 1195 2282 1196
rect 0 1143 152 1195
rect 204 1143 216 1195
rect 268 1143 280 1195
rect 332 1143 344 1195
rect 396 1143 408 1195
rect 460 1143 472 1195
rect 524 1143 536 1195
rect 588 1143 600 1195
rect 652 1143 664 1195
rect 716 1143 728 1195
rect 780 1143 792 1195
rect 844 1143 856 1195
rect 908 1143 920 1195
rect 972 1143 984 1195
rect 1036 1143 1048 1195
rect 1100 1143 1182 1195
rect 1234 1143 1246 1195
rect 1298 1143 1310 1195
rect 1362 1143 1374 1195
rect 1426 1143 1438 1195
rect 1490 1143 1502 1195
rect 1554 1143 1566 1195
rect 1618 1143 1630 1195
rect 1682 1143 1694 1195
rect 1746 1143 1758 1195
rect 1810 1143 1822 1195
rect 1874 1143 1886 1195
rect 1938 1143 1950 1195
rect 2002 1143 2014 1195
rect 2066 1143 2078 1195
rect 2130 1143 2282 1195
rect 0 1142 2282 1143
rect 0 1068 1086 1114
rect 0 1016 7 1068
rect 59 1046 1086 1068
rect 1114 1113 1168 1142
rect 1114 1061 1115 1113
rect 1167 1061 1168 1113
rect 1114 1049 1168 1061
rect 59 1016 66 1046
rect 1114 1018 1115 1049
rect 0 1004 66 1016
rect 0 952 7 1004
rect 59 962 66 1004
rect 94 997 1115 1018
rect 1167 1018 1168 1049
rect 1196 1068 2282 1114
rect 1196 1046 2223 1068
rect 1167 997 2188 1018
rect 94 990 2188 997
rect 2216 1016 2223 1046
rect 2275 1016 2282 1068
rect 2216 1004 2282 1016
rect 1114 985 1168 990
rect 59 952 1086 962
rect 0 940 1086 952
rect 0 888 7 940
rect 59 934 1086 940
rect 59 888 66 934
rect 1114 933 1115 985
rect 1167 933 1168 985
rect 2216 962 2223 1004
rect 1196 952 2223 962
rect 2275 952 2282 1004
rect 1196 940 2282 952
rect 1196 934 2223 940
rect 1114 921 1168 933
rect 1114 906 1115 921
rect 0 876 66 888
rect 94 878 1115 906
rect 0 824 7 876
rect 59 850 66 876
rect 1114 869 1115 878
rect 1167 906 1168 921
rect 1167 878 2188 906
rect 2216 888 2223 934
rect 2275 888 2282 940
rect 1167 869 1168 878
rect 1114 857 1168 869
rect 59 824 1086 850
rect 0 822 1086 824
rect 0 812 66 822
rect 0 760 7 812
rect 59 760 66 812
rect 1114 805 1115 857
rect 1167 805 1168 857
rect 2216 876 2282 888
rect 2216 850 2223 876
rect 1196 824 2223 850
rect 2275 824 2282 876
rect 1196 822 2282 824
rect 1114 794 1168 805
rect 2216 812 2282 822
rect 94 793 2188 794
rect 94 766 1115 793
rect 0 748 66 760
rect 0 696 7 748
rect 59 738 66 748
rect 1114 741 1115 766
rect 1167 766 2188 793
rect 1167 741 1168 766
rect 59 710 1086 738
rect 1114 729 1168 741
rect 2216 760 2223 812
rect 2275 760 2282 812
rect 2216 748 2282 760
rect 2216 738 2223 748
rect 59 696 66 710
rect 0 684 66 696
rect 0 632 7 684
rect 59 632 66 684
rect 1114 682 1115 729
rect 94 677 1115 682
rect 1167 682 1168 729
rect 1196 710 2223 738
rect 2216 696 2223 710
rect 2275 696 2282 748
rect 2216 684 2282 696
rect 1167 677 2188 682
rect 94 665 2188 677
rect 94 654 1115 665
rect 0 626 66 632
rect 0 620 1086 626
rect 0 568 7 620
rect 59 598 1086 620
rect 1114 613 1115 654
rect 1167 654 2188 665
rect 1167 613 1168 654
rect 2216 632 2223 684
rect 2275 632 2282 684
rect 2216 626 2282 632
rect 1114 601 1168 613
rect 59 568 66 598
rect 1114 570 1115 601
rect 0 556 66 568
rect 0 504 7 556
rect 59 514 66 556
rect 94 549 1115 570
rect 1167 570 1168 601
rect 1196 620 2282 626
rect 1196 598 2223 620
rect 1167 549 2188 570
rect 94 542 2188 549
rect 2216 568 2223 598
rect 2275 568 2282 620
rect 2216 556 2282 568
rect 1114 537 1168 542
rect 59 504 1086 514
rect 0 492 1086 504
rect 0 440 7 492
rect 59 486 1086 492
rect 59 440 66 486
rect 1114 485 1115 537
rect 1167 485 1168 537
rect 2216 514 2223 556
rect 1196 504 2223 514
rect 2275 504 2282 556
rect 1196 492 2282 504
rect 1196 486 2223 492
rect 1114 473 1168 485
rect 1114 458 1115 473
rect 0 428 66 440
rect 94 430 1115 458
rect 0 376 7 428
rect 59 402 66 428
rect 1114 421 1115 430
rect 1167 458 1168 473
rect 1167 430 2188 458
rect 2216 440 2223 486
rect 2275 440 2282 492
rect 1167 421 1168 430
rect 1114 409 1168 421
rect 59 376 1086 402
rect 0 374 1086 376
rect 0 364 66 374
rect 0 312 7 364
rect 59 312 66 364
rect 1114 357 1115 409
rect 1167 357 1168 409
rect 2216 428 2282 440
rect 2216 402 2223 428
rect 1196 376 2223 402
rect 2275 376 2282 428
rect 1196 374 2282 376
rect 1114 346 1168 357
rect 2216 364 2282 374
rect 94 345 2188 346
rect 94 318 1115 345
rect 0 300 66 312
rect 0 248 7 300
rect 59 290 66 300
rect 1114 293 1115 318
rect 1167 318 2188 345
rect 1167 293 1168 318
rect 59 262 1086 290
rect 1114 281 1168 293
rect 2216 312 2223 364
rect 2275 312 2282 364
rect 2216 300 2282 312
rect 2216 290 2223 300
rect 59 248 66 262
rect 0 236 66 248
rect 0 184 7 236
rect 59 184 66 236
rect 1114 234 1115 281
rect 94 229 1115 234
rect 1167 234 1168 281
rect 1196 262 2223 290
rect 2216 248 2223 262
rect 2275 248 2282 300
rect 2216 236 2282 248
rect 1167 229 2188 234
rect 94 217 2188 229
rect 94 206 1115 217
rect 0 178 66 184
rect 0 172 1086 178
rect 0 120 7 172
rect 59 150 1086 172
rect 1114 165 1115 206
rect 1167 206 2188 217
rect 1167 165 1168 206
rect 2216 184 2223 236
rect 2275 184 2282 236
rect 2216 178 2282 184
rect 1114 153 1168 165
rect 59 120 66 150
rect 1114 122 1115 153
rect 0 108 66 120
rect 0 56 7 108
rect 59 66 66 108
rect 94 101 1115 122
rect 1167 122 1168 153
rect 1196 172 2282 178
rect 1196 150 2223 172
rect 1167 101 2188 122
rect 94 94 2188 101
rect 2216 120 2223 150
rect 2275 120 2282 172
rect 2216 108 2282 120
rect 59 59 1086 66
rect 59 56 88 59
rect 0 7 88 56
rect 140 7 152 59
rect 204 7 216 59
rect 268 7 280 59
rect 332 7 344 59
rect 396 7 408 59
rect 460 7 472 59
rect 524 7 536 59
rect 588 7 600 59
rect 652 7 664 59
rect 716 7 728 59
rect 780 7 792 59
rect 844 7 856 59
rect 908 7 920 59
rect 972 7 984 59
rect 1036 7 1086 59
rect 0 0 1086 7
rect 1114 0 1168 94
rect 2216 66 2223 108
rect 1196 59 2223 66
rect 1196 7 1246 59
rect 1298 7 1310 59
rect 1362 7 1374 59
rect 1426 7 1438 59
rect 1490 7 1502 59
rect 1554 7 1566 59
rect 1618 7 1630 59
rect 1682 7 1694 59
rect 1746 7 1758 59
rect 1810 7 1822 59
rect 1874 7 1886 59
rect 1938 7 1950 59
rect 2002 7 2014 59
rect 2066 7 2078 59
rect 2130 7 2142 59
rect 2194 56 2223 59
rect 2275 56 2282 108
rect 2194 7 2282 56
rect 1196 0 2282 7
<< labels >>
flabel metal2 s 1018 2293 1048 2321 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 1119 2288 1161 2324 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 1176 1289 1197 1338 0 FreeSans 1600 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 748694
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 719224
string device primitive
<< end >>
