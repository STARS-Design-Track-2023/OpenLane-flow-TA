magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__hvdfm1sd2__example_55959141808243  sky130_fd_pr__hvdfm1sd2__example_55959141808243_0
timestamp 1686671242
transform 1 0 180 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808243  sky130_fd_pr__hvdfm1sd2__example_55959141808243_1
timestamp 1686671242
transform 1 0 416 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808243  sky130_fd_pr__hvdfm1sd2__example_55959141808243_2
timestamp 1686671242
transform 1 0 652 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808242  sky130_fd_pr__hvdfm1sd__example_55959141808242_0
timestamp 1686671242
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808242  sky130_fd_pr__hvdfm1sd__example_55959141808242_1
timestamp 1686671242
transform 1 0 888 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 37242638
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37240094
<< end >>
