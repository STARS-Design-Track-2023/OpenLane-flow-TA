magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 26 21 612 203
rect 29 -17 63 21
<< scnmos >>
rect 108 47 138 177
rect 192 47 222 177
rect 276 47 306 177
rect 428 47 458 177
rect 500 47 530 177
<< scpmoshvt >>
rect 108 297 138 497
rect 192 297 222 497
rect 276 297 306 497
rect 396 297 426 497
rect 500 297 530 497
<< ndiff >>
rect 52 157 108 177
rect 52 123 64 157
rect 98 123 108 157
rect 52 89 108 123
rect 52 55 64 89
rect 98 55 108 89
rect 52 47 108 55
rect 138 126 192 177
rect 138 92 148 126
rect 182 92 192 126
rect 138 47 192 92
rect 222 89 276 177
rect 222 55 232 89
rect 266 55 276 89
rect 222 47 276 55
rect 306 126 428 177
rect 306 92 316 126
rect 350 92 428 126
rect 306 47 428 92
rect 458 47 500 177
rect 530 157 586 177
rect 530 123 540 157
rect 574 123 586 157
rect 530 89 586 123
rect 530 55 540 89
rect 574 55 586 89
rect 530 47 586 55
<< pdiff >>
rect 52 477 108 497
rect 52 443 64 477
rect 98 443 108 477
rect 52 409 108 443
rect 52 375 64 409
rect 98 375 108 409
rect 52 341 108 375
rect 52 307 64 341
rect 98 307 108 341
rect 52 297 108 307
rect 138 297 192 497
rect 222 297 276 497
rect 306 477 396 497
rect 306 443 334 477
rect 368 443 396 477
rect 306 409 396 443
rect 306 375 334 409
rect 368 375 396 409
rect 306 341 396 375
rect 306 307 334 341
rect 368 307 396 341
rect 306 297 396 307
rect 426 477 500 497
rect 426 443 446 477
rect 480 443 500 477
rect 426 409 500 443
rect 426 375 446 409
rect 480 375 500 409
rect 426 297 500 375
rect 530 477 592 497
rect 530 443 546 477
rect 580 443 592 477
rect 530 409 592 443
rect 530 375 546 409
rect 580 375 592 409
rect 530 341 592 375
rect 530 307 546 341
rect 580 307 592 341
rect 530 297 592 307
<< ndiffc >>
rect 64 123 98 157
rect 64 55 98 89
rect 148 92 182 126
rect 232 55 266 89
rect 316 92 350 126
rect 540 123 574 157
rect 540 55 574 89
<< pdiffc >>
rect 64 443 98 477
rect 64 375 98 409
rect 64 307 98 341
rect 334 443 368 477
rect 334 375 368 409
rect 334 307 368 341
rect 446 443 480 477
rect 446 375 480 409
rect 546 443 580 477
rect 546 375 580 409
rect 546 307 580 341
<< poly >>
rect 108 497 138 523
rect 192 497 222 523
rect 276 497 306 523
rect 396 497 426 523
rect 500 497 530 523
rect 108 265 138 297
rect 192 265 222 297
rect 276 265 306 297
rect 396 265 426 297
rect 500 265 530 297
rect 54 249 138 265
rect 54 215 64 249
rect 98 215 138 249
rect 54 199 138 215
rect 180 249 234 265
rect 180 215 190 249
rect 224 215 234 249
rect 180 199 234 215
rect 276 249 330 265
rect 276 215 286 249
rect 320 215 330 249
rect 276 199 330 215
rect 396 249 458 265
rect 396 215 406 249
rect 440 215 458 249
rect 396 199 458 215
rect 108 177 138 199
rect 192 177 222 199
rect 276 177 306 199
rect 428 177 458 199
rect 500 249 610 265
rect 500 215 566 249
rect 600 215 610 249
rect 500 199 610 215
rect 500 177 530 199
rect 108 21 138 47
rect 192 21 222 47
rect 276 21 306 47
rect 428 21 458 47
rect 500 21 530 47
<< polycont >>
rect 64 215 98 249
rect 190 215 224 249
rect 286 215 320 249
rect 406 215 440 249
rect 566 215 600 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 477 156 527
rect 17 443 64 477
rect 98 443 156 477
rect 17 409 156 443
rect 17 375 64 409
rect 98 375 156 409
rect 17 341 156 375
rect 17 307 64 341
rect 98 307 156 341
rect 17 299 156 307
rect 17 249 156 265
rect 17 215 64 249
rect 98 215 156 249
rect 17 199 156 215
rect 190 249 252 493
rect 286 477 396 493
rect 286 443 334 477
rect 368 443 396 477
rect 286 409 396 443
rect 286 375 334 409
rect 368 375 396 409
rect 286 341 396 375
rect 430 477 496 527
rect 430 443 446 477
rect 480 443 496 477
rect 430 409 496 443
rect 430 375 446 409
rect 480 375 496 409
rect 430 367 496 375
rect 530 477 627 493
rect 530 443 546 477
rect 580 443 627 477
rect 530 409 627 443
rect 530 375 546 409
rect 580 375 627 409
rect 286 307 334 341
rect 368 333 396 341
rect 530 341 627 375
rect 530 333 546 341
rect 368 307 546 333
rect 580 307 627 341
rect 286 299 627 307
rect 224 215 252 249
rect 190 199 252 215
rect 286 249 356 265
rect 320 215 356 249
rect 286 199 356 215
rect 397 249 440 265
rect 397 215 406 249
rect 17 157 114 165
rect 17 123 64 157
rect 98 123 114 157
rect 17 89 114 123
rect 17 55 64 89
rect 98 55 114 89
rect 17 17 114 55
rect 148 131 350 165
rect 148 126 182 131
rect 316 126 350 131
rect 148 51 182 92
rect 216 89 282 97
rect 216 55 232 89
rect 266 55 282 89
rect 216 17 282 55
rect 316 51 350 92
rect 397 64 440 215
rect 489 165 532 299
rect 566 249 627 265
rect 600 215 627 249
rect 566 199 627 215
rect 489 157 627 165
rect 489 123 540 157
rect 574 123 627 157
rect 489 89 627 123
rect 489 55 540 89
rect 574 55 627 89
rect 489 51 627 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 581 85 615 119 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 489 153 523 187 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 489 85 523 119 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 489 289 523 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 305 357 339 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 305 425 339 459 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 581 425 615 459 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 581 357 615 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o311ai_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 884638
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 877790
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.220 0.000 
<< end >>
