magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1103 203
rect 30 -17 64 21
<< locali >>
rect 86 199 148 265
rect 296 199 350 323
rect 393 199 487 265
rect 536 199 679 265
rect 783 349 817 493
rect 951 349 985 493
rect 783 315 1086 349
rect 114 161 148 199
rect 536 161 570 199
rect 114 127 570 161
rect 1040 161 1086 315
rect 783 127 1086 161
rect 783 51 817 127
rect 951 51 985 127
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 18 333 69 493
rect 103 367 164 527
rect 198 455 554 489
rect 198 387 268 455
rect 615 421 649 493
rect 683 451 749 527
rect 306 387 649 421
rect 713 353 747 357
rect 18 299 216 333
rect 18 125 52 299
rect 182 199 216 299
rect 396 319 747 353
rect 713 249 747 319
rect 851 383 917 527
rect 1019 383 1085 527
rect 713 215 1006 249
rect 713 165 747 215
rect 612 131 747 165
rect 18 59 69 125
rect 612 93 646 131
rect 103 17 169 93
rect 395 59 646 93
rect 683 17 749 93
rect 851 17 917 93
rect 1019 17 1085 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 296 199 350 323 6 A0
port 1 nsew signal input
rlabel locali s 393 199 487 265 6 A1
port 2 nsew signal input
rlabel locali s 114 127 570 161 6 S
port 3 nsew signal input
rlabel locali s 536 161 570 199 6 S
port 3 nsew signal input
rlabel locali s 536 199 679 265 6 S
port 3 nsew signal input
rlabel locali s 114 161 148 199 6 S
port 3 nsew signal input
rlabel locali s 86 199 148 265 6 S
port 3 nsew signal input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1103 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 951 51 985 127 6 X
port 8 nsew signal output
rlabel locali s 783 51 817 127 6 X
port 8 nsew signal output
rlabel locali s 783 127 1086 161 6 X
port 8 nsew signal output
rlabel locali s 1040 161 1086 315 6 X
port 8 nsew signal output
rlabel locali s 783 315 1086 349 6 X
port 8 nsew signal output
rlabel locali s 951 349 985 493 6 X
port 8 nsew signal output
rlabel locali s 783 349 817 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1690600
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1682266
<< end >>
