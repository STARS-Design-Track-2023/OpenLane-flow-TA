magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 4 21 367 203
rect 29 -17 63 21
<< scnmos >>
rect 83 47 113 177
rect 169 47 199 177
rect 258 47 288 177
<< scpmoshvt >>
rect 83 297 113 497
rect 169 297 199 497
rect 258 297 288 497
<< ndiff >>
rect 30 93 83 177
rect 30 59 38 93
rect 72 59 83 93
rect 30 47 83 59
rect 113 127 169 177
rect 113 93 124 127
rect 158 93 169 127
rect 113 47 169 93
rect 199 47 258 177
rect 288 123 341 177
rect 288 89 299 123
rect 333 89 341 123
rect 288 47 341 89
<< pdiff >>
rect 30 453 83 497
rect 30 419 38 453
rect 72 419 83 453
rect 30 379 83 419
rect 30 345 38 379
rect 72 345 83 379
rect 30 297 83 345
rect 113 475 169 497
rect 113 441 124 475
rect 158 441 169 475
rect 113 407 169 441
rect 113 373 124 407
rect 158 373 169 407
rect 113 297 169 373
rect 199 489 258 497
rect 199 455 210 489
rect 244 455 258 489
rect 199 297 258 455
rect 288 483 341 497
rect 288 449 299 483
rect 333 449 341 483
rect 288 415 341 449
rect 288 381 299 415
rect 333 381 341 415
rect 288 347 341 381
rect 288 313 299 347
rect 333 313 341 347
rect 288 297 341 313
<< ndiffc >>
rect 38 59 72 93
rect 124 93 158 127
rect 299 89 333 123
<< pdiffc >>
rect 38 419 72 453
rect 38 345 72 379
rect 124 441 158 475
rect 124 373 158 407
rect 210 455 244 489
rect 299 449 333 483
rect 299 381 333 415
rect 299 313 333 347
<< poly >>
rect 83 497 113 523
rect 169 497 199 523
rect 258 497 288 523
rect 83 265 113 297
rect 169 265 199 297
rect 258 265 288 297
rect 21 249 113 265
rect 21 215 31 249
rect 65 215 113 249
rect 21 199 113 215
rect 162 249 216 265
rect 162 215 172 249
rect 206 215 216 249
rect 162 199 216 215
rect 258 249 342 265
rect 258 215 298 249
rect 332 215 342 249
rect 258 199 342 215
rect 83 177 113 199
rect 169 177 199 199
rect 258 177 288 199
rect 83 21 113 47
rect 169 21 199 47
rect 258 21 288 47
<< polycont >>
rect 31 215 65 249
rect 172 215 206 249
rect 298 215 332 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 19 453 74 491
rect 19 419 38 453
rect 72 419 74 453
rect 19 379 74 419
rect 19 345 38 379
rect 72 345 74 379
rect 108 475 174 491
rect 108 441 124 475
rect 158 441 174 475
rect 108 407 174 441
rect 208 489 247 527
rect 208 455 210 489
rect 244 455 247 489
rect 208 439 247 455
rect 283 483 349 491
rect 283 449 299 483
rect 333 449 349 483
rect 108 373 124 407
rect 158 405 174 407
rect 283 415 349 449
rect 283 405 299 415
rect 158 381 299 405
rect 333 381 349 415
rect 158 373 349 381
rect 108 371 349 373
rect 19 337 74 345
rect 170 347 349 371
rect 19 299 136 337
rect 170 313 299 347
rect 333 313 349 347
rect 170 305 349 313
rect 19 249 67 265
rect 19 215 31 249
rect 65 215 67 249
rect 19 135 67 215
rect 101 165 136 299
rect 170 249 253 265
rect 170 215 172 249
rect 206 215 253 249
rect 170 199 253 215
rect 289 249 348 265
rect 289 215 298 249
rect 332 215 348 249
rect 289 199 348 215
rect 101 129 167 165
rect 122 127 167 129
rect 22 93 88 95
rect 22 59 38 93
rect 72 59 88 93
rect 22 17 88 59
rect 122 93 124 127
rect 158 93 167 127
rect 122 53 167 93
rect 207 75 253 199
rect 289 123 349 163
rect 289 89 299 123
rect 333 89 349 123
rect 289 17 349 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 213 153 247 187 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 213 85 247 119 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 29 425 63 459 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 29 357 63 391 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a21oi_1
rlabel metal1 s 0 -48 368 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 368 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_END 4042676
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4038006
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 9.200 13.600 
<< end >>
