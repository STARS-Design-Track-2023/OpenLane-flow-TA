magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect 2009 2487 2390 3309
rect 1423 1767 2661 1843
rect -216 1759 2661 1767
rect -216 1388 5375 1759
rect -216 1214 5268 1388
rect -251 521 5268 1214
rect -251 513 2628 521
rect 1316 440 2628 513
<< pwell >>
rect 2069 3651 2337 3737
rect 2072 3606 2337 3651
rect 2072 3414 2350 3606
rect 2758 2205 3740 2311
rect 1463 2172 3740 2205
rect 280 2164 3740 2172
rect 280 2086 5196 2164
rect 280 2064 1285 2086
rect -176 1872 1285 2064
rect 1463 2013 5196 2086
rect 2783 1864 5196 2013
rect -176 216 1230 408
rect 291 177 1230 216
rect 1430 177 2588 270
rect 2783 202 5193 416
rect 291 91 2588 177
rect 2779 116 5193 202
rect 1430 78 2588 91
<< mvnmos >>
rect 2151 3440 2271 3580
rect 1542 2039 1662 2179
rect 1718 2039 1838 2179
rect 1894 2039 2014 2179
rect 2070 2039 2190 2179
rect 2246 2039 2366 2179
rect 2422 2039 2542 2179
rect -97 1898 23 2038
rect 79 1898 199 2038
rect 379 1898 499 2038
rect 555 1898 675 2038
rect 731 1898 851 2038
rect 907 1898 1027 2038
rect 1083 1898 1203 2038
rect 2862 1890 2982 2030
rect 3038 1890 3158 2030
rect 3214 1890 3334 2030
rect 3514 1890 3634 2030
rect 3690 1890 3810 2030
rect 3866 1890 3986 2030
rect 4042 1890 4162 2030
rect 4342 1890 4462 2030
rect 4518 1890 4638 2030
rect 4818 1890 4938 2030
rect 4994 1890 5114 2030
rect -97 242 23 382
rect 79 242 199 382
rect 379 242 499 382
rect 555 242 675 382
rect 731 242 851 382
rect 1031 242 1151 382
rect 2862 250 2982 390
rect 3038 250 3158 390
rect 3214 250 3334 390
rect 3514 250 3634 390
rect 3690 250 3810 390
rect 3990 250 4110 390
rect 4166 250 4286 390
rect 4342 250 4462 390
rect 4518 250 4638 390
rect 4818 250 4938 390
rect 4994 250 5114 390
rect 1509 104 1629 244
rect 1685 104 1805 244
rect 1861 104 1981 244
rect 2037 104 2157 244
rect 2213 104 2333 244
rect 2389 104 2509 244
<< mvpmos >>
rect 2151 3042 2271 3242
rect 2151 2774 2271 2974
rect -97 1500 23 1700
rect 79 1500 199 1700
rect 379 1500 499 1700
rect 555 1500 675 1700
rect 731 1500 851 1700
rect 907 1500 1027 1700
rect 1083 1500 1203 1700
rect 1542 1577 1662 1777
rect 1718 1577 1838 1777
rect 1894 1577 2014 1777
rect 2070 1577 2190 1777
rect 2246 1577 2366 1777
rect 2422 1577 2542 1777
rect -97 1232 23 1432
rect 79 1232 199 1432
rect 379 1232 499 1432
rect 555 1232 675 1432
rect 731 1232 851 1432
rect 907 1232 1027 1432
rect 1083 1232 1203 1432
rect 1542 1309 1662 1509
rect 1718 1309 1838 1509
rect 1894 1309 2014 1509
rect 2070 1309 2190 1509
rect 2246 1309 2366 1509
rect 2422 1309 2542 1509
rect 2862 1492 2982 1692
rect 3038 1492 3158 1692
rect 3214 1492 3334 1692
rect 3514 1492 3634 1692
rect 3690 1492 3810 1692
rect 3866 1492 3986 1692
rect 4042 1492 4162 1692
rect 4342 1492 4462 1692
rect 4518 1492 4638 1692
rect 4818 1492 4938 1692
rect 4994 1492 5114 1692
rect 2862 1224 2982 1424
rect 3038 1224 3158 1424
rect 3214 1224 3334 1424
rect 3514 1224 3634 1424
rect 3690 1224 3810 1424
rect 3866 1224 3986 1424
rect 4042 1224 4162 1424
rect 4342 1224 4462 1424
rect 4518 1224 4638 1424
rect 4818 1224 4938 1424
rect 4994 1224 5114 1424
rect -97 848 23 1048
rect 79 848 199 1048
rect 379 848 499 1048
rect 555 848 675 1048
rect 731 848 851 1048
rect 1031 848 1151 1048
rect -97 580 23 780
rect 79 580 199 780
rect 379 580 499 780
rect 555 580 675 780
rect 731 580 851 780
rect 1031 580 1151 780
rect 1509 774 1629 974
rect 1685 774 1805 974
rect 1861 774 1981 974
rect 2037 774 2157 974
rect 2213 774 2333 974
rect 2389 774 2509 974
rect 2862 856 2982 1056
rect 3038 856 3158 1056
rect 3214 856 3334 1056
rect 3514 856 3634 1056
rect 3690 856 3810 1056
rect 3990 856 4110 1056
rect 4166 856 4286 1056
rect 4342 856 4462 1056
rect 4518 856 4638 1056
rect 4818 856 4938 1056
rect 4994 856 5114 1056
rect 1509 506 1629 706
rect 1685 506 1805 706
rect 1861 506 1981 706
rect 2037 506 2157 706
rect 2213 506 2333 706
rect 2389 506 2509 706
rect 2862 588 2982 788
rect 3038 588 3158 788
rect 3214 588 3334 788
rect 3514 588 3634 788
rect 3690 588 3810 788
rect 3990 588 4110 788
rect 4166 588 4286 788
rect 4342 588 4462 788
rect 4518 588 4638 788
rect 4818 588 4938 788
rect 4994 588 5114 788
<< mvndiff >>
rect 2098 3554 2151 3580
rect 2098 3520 2106 3554
rect 2140 3520 2151 3554
rect 2098 3486 2151 3520
rect 2098 3452 2106 3486
rect 2140 3452 2151 3486
rect 2098 3440 2151 3452
rect 2271 3554 2324 3580
rect 2271 3520 2282 3554
rect 2316 3520 2324 3554
rect 2271 3486 2324 3520
rect 2271 3452 2282 3486
rect 2316 3452 2324 3486
rect 2271 3440 2324 3452
rect 1489 2167 1542 2179
rect 1489 2133 1497 2167
rect 1531 2133 1542 2167
rect 1489 2099 1542 2133
rect 1489 2065 1497 2099
rect 1531 2065 1542 2099
rect 1489 2039 1542 2065
rect 1662 2167 1718 2179
rect 1662 2133 1673 2167
rect 1707 2133 1718 2167
rect 1662 2099 1718 2133
rect 1662 2065 1673 2099
rect 1707 2065 1718 2099
rect 1662 2039 1718 2065
rect 1838 2167 1894 2179
rect 1838 2133 1849 2167
rect 1883 2133 1894 2167
rect 1838 2099 1894 2133
rect 1838 2065 1849 2099
rect 1883 2065 1894 2099
rect 1838 2039 1894 2065
rect 2014 2167 2070 2179
rect 2014 2133 2025 2167
rect 2059 2133 2070 2167
rect 2014 2099 2070 2133
rect 2014 2065 2025 2099
rect 2059 2065 2070 2099
rect 2014 2039 2070 2065
rect 2190 2167 2246 2179
rect 2190 2133 2201 2167
rect 2235 2133 2246 2167
rect 2190 2099 2246 2133
rect 2190 2065 2201 2099
rect 2235 2065 2246 2099
rect 2190 2039 2246 2065
rect 2366 2167 2422 2179
rect 2366 2133 2377 2167
rect 2411 2133 2422 2167
rect 2366 2099 2422 2133
rect 2366 2065 2377 2099
rect 2411 2065 2422 2099
rect 2366 2039 2422 2065
rect 2542 2167 2595 2179
rect 2542 2133 2553 2167
rect 2587 2133 2595 2167
rect 2542 2099 2595 2133
rect 2542 2065 2553 2099
rect 2587 2065 2595 2099
rect 2542 2039 2595 2065
rect -150 2012 -97 2038
rect -150 1978 -142 2012
rect -108 1978 -97 2012
rect -150 1944 -97 1978
rect -150 1910 -142 1944
rect -108 1910 -97 1944
rect -150 1898 -97 1910
rect 23 2012 79 2038
rect 23 1978 34 2012
rect 68 1978 79 2012
rect 23 1944 79 1978
rect 23 1910 34 1944
rect 68 1910 79 1944
rect 23 1898 79 1910
rect 199 2012 255 2038
rect 199 1978 210 2012
rect 244 1978 255 2012
rect 199 1944 255 1978
rect 199 1910 210 1944
rect 244 1910 255 1944
rect 199 1898 255 1910
rect 326 2012 379 2038
rect 326 1978 334 2012
rect 368 1978 379 2012
rect 326 1944 379 1978
rect 326 1910 334 1944
rect 368 1910 379 1944
rect 326 1898 379 1910
rect 499 2012 555 2038
rect 499 1978 510 2012
rect 544 1978 555 2012
rect 499 1944 555 1978
rect 499 1910 510 1944
rect 544 1910 555 1944
rect 499 1898 555 1910
rect 675 2012 731 2038
rect 675 1978 686 2012
rect 720 1978 731 2012
rect 675 1944 731 1978
rect 675 1910 686 1944
rect 720 1910 731 1944
rect 675 1898 731 1910
rect 851 2012 907 2038
rect 851 1978 862 2012
rect 896 1978 907 2012
rect 851 1944 907 1978
rect 851 1910 862 1944
rect 896 1910 907 1944
rect 851 1898 907 1910
rect 1027 2012 1083 2038
rect 1027 1978 1038 2012
rect 1072 1978 1083 2012
rect 1027 1944 1083 1978
rect 1027 1910 1038 1944
rect 1072 1910 1083 1944
rect 1027 1898 1083 1910
rect 1203 2012 1259 2038
rect 1203 1978 1214 2012
rect 1248 1978 1259 2012
rect 1203 1944 1259 1978
rect 1203 1910 1214 1944
rect 1248 1910 1259 1944
rect 1203 1898 1259 1910
rect 2809 2004 2862 2030
rect 2809 1970 2817 2004
rect 2851 1970 2862 2004
rect 2809 1936 2862 1970
rect 2809 1902 2817 1936
rect 2851 1902 2862 1936
rect 2809 1890 2862 1902
rect 2982 2004 3038 2030
rect 2982 1970 2993 2004
rect 3027 1970 3038 2004
rect 2982 1936 3038 1970
rect 2982 1902 2993 1936
rect 3027 1902 3038 1936
rect 2982 1890 3038 1902
rect 3158 2004 3214 2030
rect 3158 1970 3169 2004
rect 3203 1970 3214 2004
rect 3158 1936 3214 1970
rect 3158 1902 3169 1936
rect 3203 1902 3214 1936
rect 3158 1890 3214 1902
rect 3334 2004 3387 2030
rect 3334 1970 3345 2004
rect 3379 1970 3387 2004
rect 3334 1936 3387 1970
rect 3334 1902 3345 1936
rect 3379 1902 3387 1936
rect 3334 1890 3387 1902
rect 3461 2004 3514 2030
rect 3461 1970 3469 2004
rect 3503 1970 3514 2004
rect 3461 1936 3514 1970
rect 3461 1902 3469 1936
rect 3503 1902 3514 1936
rect 3461 1890 3514 1902
rect 3634 1890 3690 2030
rect 3810 2004 3866 2030
rect 3810 1970 3821 2004
rect 3855 1970 3866 2004
rect 3810 1936 3866 1970
rect 3810 1902 3821 1936
rect 3855 1902 3866 1936
rect 3810 1890 3866 1902
rect 3986 1890 4042 2030
rect 4162 2004 4215 2030
rect 4162 1970 4173 2004
rect 4207 1970 4215 2004
rect 4162 1936 4215 1970
rect 4162 1902 4173 1936
rect 4207 1902 4215 1936
rect 4162 1890 4215 1902
rect 4289 2004 4342 2030
rect 4289 1970 4297 2004
rect 4331 1970 4342 2004
rect 4289 1936 4342 1970
rect 4289 1902 4297 1936
rect 4331 1902 4342 1936
rect 4289 1890 4342 1902
rect 4462 1890 4518 2030
rect 4638 2004 4691 2030
rect 4638 1970 4649 2004
rect 4683 1970 4691 2004
rect 4638 1936 4691 1970
rect 4638 1902 4649 1936
rect 4683 1902 4691 1936
rect 4638 1890 4691 1902
rect 4765 2004 4818 2030
rect 4765 1970 4773 2004
rect 4807 1970 4818 2004
rect 4765 1936 4818 1970
rect 4765 1902 4773 1936
rect 4807 1902 4818 1936
rect 4765 1890 4818 1902
rect 4938 2004 4994 2030
rect 4938 1970 4949 2004
rect 4983 1970 4994 2004
rect 4938 1936 4994 1970
rect 4938 1902 4949 1936
rect 4983 1902 4994 1936
rect 4938 1890 4994 1902
rect 5114 2004 5170 2030
rect 5114 1970 5125 2004
rect 5159 1970 5170 2004
rect 5114 1936 5170 1970
rect 5114 1902 5125 1936
rect 5159 1902 5170 1936
rect 5114 1890 5170 1902
rect -150 370 -97 382
rect -150 336 -142 370
rect -108 336 -97 370
rect -150 302 -97 336
rect -150 268 -142 302
rect -108 268 -97 302
rect -150 242 -97 268
rect 23 242 79 382
rect 199 370 252 382
rect 199 336 210 370
rect 244 336 252 370
rect 199 302 252 336
rect 199 268 210 302
rect 244 268 252 302
rect 199 242 252 268
rect 326 370 379 382
rect 326 336 334 370
rect 368 336 379 370
rect 326 302 379 336
rect 326 268 334 302
rect 368 268 379 302
rect 326 242 379 268
rect 499 370 555 382
rect 499 336 510 370
rect 544 336 555 370
rect 499 302 555 336
rect 499 268 510 302
rect 544 268 555 302
rect 499 242 555 268
rect 675 370 731 382
rect 675 336 686 370
rect 720 336 731 370
rect 675 302 731 336
rect 675 268 686 302
rect 720 268 731 302
rect 675 242 731 268
rect 851 370 904 382
rect 851 336 862 370
rect 896 336 904 370
rect 851 302 904 336
rect 851 268 862 302
rect 896 268 904 302
rect 851 242 904 268
rect 978 370 1031 382
rect 978 336 986 370
rect 1020 336 1031 370
rect 978 302 1031 336
rect 978 268 986 302
rect 1020 268 1031 302
rect 978 242 1031 268
rect 1151 370 1204 382
rect 1151 336 1162 370
rect 1196 336 1204 370
rect 1151 302 1204 336
rect 1151 268 1162 302
rect 1196 268 1204 302
rect 1151 242 1204 268
rect 2809 378 2862 390
rect 2809 344 2817 378
rect 2851 344 2862 378
rect 2809 310 2862 344
rect 2809 276 2817 310
rect 2851 276 2862 310
rect 2809 250 2862 276
rect 2982 378 3038 390
rect 2982 344 2993 378
rect 3027 344 3038 378
rect 2982 310 3038 344
rect 2982 276 2993 310
rect 3027 276 3038 310
rect 2982 250 3038 276
rect 3158 378 3214 390
rect 3158 344 3169 378
rect 3203 344 3214 378
rect 3158 310 3214 344
rect 3158 276 3169 310
rect 3203 276 3214 310
rect 3158 250 3214 276
rect 3334 378 3387 390
rect 3334 344 3345 378
rect 3379 344 3387 378
rect 3334 310 3387 344
rect 3334 276 3345 310
rect 3379 276 3387 310
rect 3334 250 3387 276
rect 3461 378 3514 390
rect 3461 344 3469 378
rect 3503 344 3514 378
rect 3461 310 3514 344
rect 3461 276 3469 310
rect 3503 276 3514 310
rect 3461 250 3514 276
rect 3634 250 3690 390
rect 3810 378 3863 390
rect 3810 344 3821 378
rect 3855 344 3863 378
rect 3810 310 3863 344
rect 3810 276 3821 310
rect 3855 276 3863 310
rect 3810 250 3863 276
rect 3937 378 3990 390
rect 3937 344 3945 378
rect 3979 344 3990 378
rect 3937 310 3990 344
rect 3937 276 3945 310
rect 3979 276 3990 310
rect 3937 250 3990 276
rect 4110 250 4166 390
rect 4286 378 4342 390
rect 4286 344 4297 378
rect 4331 344 4342 378
rect 4286 310 4342 344
rect 4286 276 4297 310
rect 4331 276 4342 310
rect 4286 250 4342 276
rect 4462 250 4518 390
rect 4638 378 4691 390
rect 4638 344 4649 378
rect 4683 344 4691 378
rect 4638 310 4691 344
rect 4638 276 4649 310
rect 4683 276 4691 310
rect 4638 250 4691 276
rect 4765 378 4818 390
rect 4765 344 4773 378
rect 4807 344 4818 378
rect 4765 310 4818 344
rect 4765 276 4773 310
rect 4807 276 4818 310
rect 4765 250 4818 276
rect 4938 250 4994 390
rect 5114 378 5167 390
rect 5114 344 5125 378
rect 5159 344 5167 378
rect 5114 310 5167 344
rect 5114 276 5125 310
rect 5159 276 5167 310
rect 5114 250 5167 276
rect 1456 218 1509 244
rect 1456 184 1464 218
rect 1498 184 1509 218
rect 1456 150 1509 184
rect 1456 116 1464 150
rect 1498 116 1509 150
rect 1456 104 1509 116
rect 1629 218 1685 244
rect 1629 184 1640 218
rect 1674 184 1685 218
rect 1629 150 1685 184
rect 1629 116 1640 150
rect 1674 116 1685 150
rect 1629 104 1685 116
rect 1805 218 1861 244
rect 1805 184 1816 218
rect 1850 184 1861 218
rect 1805 150 1861 184
rect 1805 116 1816 150
rect 1850 116 1861 150
rect 1805 104 1861 116
rect 1981 218 2037 244
rect 1981 184 1992 218
rect 2026 184 2037 218
rect 1981 150 2037 184
rect 1981 116 1992 150
rect 2026 116 2037 150
rect 1981 104 2037 116
rect 2157 218 2213 244
rect 2157 184 2168 218
rect 2202 184 2213 218
rect 2157 150 2213 184
rect 2157 116 2168 150
rect 2202 116 2213 150
rect 2157 104 2213 116
rect 2333 218 2389 244
rect 2333 184 2344 218
rect 2378 184 2389 218
rect 2333 150 2389 184
rect 2333 116 2344 150
rect 2378 116 2389 150
rect 2333 104 2389 116
rect 2509 218 2562 244
rect 2509 184 2520 218
rect 2554 184 2562 218
rect 2509 150 2562 184
rect 2509 116 2520 150
rect 2554 116 2562 150
rect 2509 104 2562 116
<< mvpdiff >>
rect 2098 3224 2151 3242
rect 2098 3190 2106 3224
rect 2140 3190 2151 3224
rect 2098 3156 2151 3190
rect 2098 3122 2106 3156
rect 2140 3122 2151 3156
rect 2098 3088 2151 3122
rect 2098 3054 2106 3088
rect 2140 3054 2151 3088
rect 2098 3042 2151 3054
rect 2271 3224 2324 3242
rect 2271 3190 2282 3224
rect 2316 3190 2324 3224
rect 2271 3156 2324 3190
rect 2271 3122 2282 3156
rect 2316 3122 2324 3156
rect 2271 3088 2324 3122
rect 2271 3054 2282 3088
rect 2316 3054 2324 3088
rect 2271 3042 2324 3054
rect 2098 2962 2151 2974
rect 2098 2928 2106 2962
rect 2140 2928 2151 2962
rect 2098 2894 2151 2928
rect 2098 2860 2106 2894
rect 2140 2860 2151 2894
rect 2098 2826 2151 2860
rect 2098 2792 2106 2826
rect 2140 2792 2151 2826
rect 2098 2774 2151 2792
rect 2271 2962 2324 2974
rect 2271 2928 2282 2962
rect 2316 2928 2324 2962
rect 2271 2894 2324 2928
rect 2271 2860 2282 2894
rect 2316 2860 2324 2894
rect 2271 2826 2324 2860
rect 2271 2792 2282 2826
rect 2316 2792 2324 2826
rect 2271 2774 2324 2792
rect 1489 1765 1542 1777
rect 1489 1731 1497 1765
rect 1531 1731 1542 1765
rect -150 1682 -97 1700
rect -150 1648 -142 1682
rect -108 1648 -97 1682
rect -150 1614 -97 1648
rect -150 1580 -142 1614
rect -108 1580 -97 1614
rect -150 1546 -97 1580
rect -150 1512 -142 1546
rect -108 1512 -97 1546
rect -150 1500 -97 1512
rect 23 1614 79 1700
rect 23 1580 34 1614
rect 68 1580 79 1614
rect 23 1546 79 1580
rect 23 1512 34 1546
rect 68 1512 79 1546
rect 23 1500 79 1512
rect 199 1682 252 1700
rect 199 1648 210 1682
rect 244 1648 252 1682
rect 199 1614 252 1648
rect 199 1580 210 1614
rect 244 1580 252 1614
rect 199 1546 252 1580
rect 199 1512 210 1546
rect 244 1512 252 1546
rect 199 1500 252 1512
rect 326 1682 379 1700
rect 326 1648 334 1682
rect 368 1648 379 1682
rect 326 1614 379 1648
rect 326 1580 334 1614
rect 368 1580 379 1614
rect 326 1546 379 1580
rect 326 1512 334 1546
rect 368 1512 379 1546
rect 326 1500 379 1512
rect 499 1682 555 1700
rect 499 1648 510 1682
rect 544 1648 555 1682
rect 499 1614 555 1648
rect 499 1580 510 1614
rect 544 1580 555 1614
rect 499 1546 555 1580
rect 499 1512 510 1546
rect 544 1512 555 1546
rect 499 1500 555 1512
rect 675 1682 731 1700
rect 675 1648 686 1682
rect 720 1648 731 1682
rect 675 1614 731 1648
rect 675 1580 686 1614
rect 720 1580 731 1614
rect 675 1546 731 1580
rect 675 1512 686 1546
rect 720 1512 731 1546
rect 675 1500 731 1512
rect 851 1682 907 1700
rect 851 1648 862 1682
rect 896 1648 907 1682
rect 851 1614 907 1648
rect 851 1580 862 1614
rect 896 1580 907 1614
rect 851 1546 907 1580
rect 851 1512 862 1546
rect 896 1512 907 1546
rect 851 1500 907 1512
rect 1027 1614 1083 1700
rect 1027 1580 1038 1614
rect 1072 1580 1083 1614
rect 1027 1546 1083 1580
rect 1027 1512 1038 1546
rect 1072 1512 1083 1546
rect 1027 1500 1083 1512
rect 1203 1682 1256 1700
rect 1203 1648 1214 1682
rect 1248 1648 1256 1682
rect 1203 1614 1256 1648
rect 1203 1580 1214 1614
rect 1248 1580 1256 1614
rect 1203 1546 1256 1580
rect 1489 1697 1542 1731
rect 1489 1663 1497 1697
rect 1531 1663 1542 1697
rect 1489 1629 1542 1663
rect 1489 1595 1497 1629
rect 1531 1595 1542 1629
rect 1489 1577 1542 1595
rect 1662 1765 1718 1777
rect 1662 1731 1673 1765
rect 1707 1731 1718 1765
rect 1662 1697 1718 1731
rect 1662 1663 1673 1697
rect 1707 1663 1718 1697
rect 1662 1629 1718 1663
rect 1662 1595 1673 1629
rect 1707 1595 1718 1629
rect 1662 1577 1718 1595
rect 1838 1765 1894 1777
rect 1838 1731 1849 1765
rect 1883 1731 1894 1765
rect 1838 1697 1894 1731
rect 1838 1663 1849 1697
rect 1883 1663 1894 1697
rect 1838 1629 1894 1663
rect 1838 1595 1849 1629
rect 1883 1595 1894 1629
rect 1838 1577 1894 1595
rect 2014 1765 2070 1777
rect 2014 1731 2025 1765
rect 2059 1731 2070 1765
rect 2014 1697 2070 1731
rect 2014 1663 2025 1697
rect 2059 1663 2070 1697
rect 2014 1629 2070 1663
rect 2014 1595 2025 1629
rect 2059 1595 2070 1629
rect 2014 1577 2070 1595
rect 2190 1765 2246 1777
rect 2190 1731 2201 1765
rect 2235 1731 2246 1765
rect 2190 1697 2246 1731
rect 2190 1663 2201 1697
rect 2235 1663 2246 1697
rect 2190 1629 2246 1663
rect 2190 1595 2201 1629
rect 2235 1595 2246 1629
rect 2190 1577 2246 1595
rect 2366 1765 2422 1777
rect 2366 1731 2377 1765
rect 2411 1731 2422 1765
rect 2366 1697 2422 1731
rect 2366 1663 2377 1697
rect 2411 1663 2422 1697
rect 2366 1629 2422 1663
rect 2366 1595 2377 1629
rect 2411 1595 2422 1629
rect 2366 1577 2422 1595
rect 2542 1765 2595 1777
rect 2542 1731 2553 1765
rect 2587 1731 2595 1765
rect 2542 1697 2595 1731
rect 2542 1663 2553 1697
rect 2587 1663 2595 1697
rect 2542 1629 2595 1663
rect 2542 1595 2553 1629
rect 2587 1595 2595 1629
rect 2542 1577 2595 1595
rect 2809 1674 2862 1692
rect 2809 1640 2817 1674
rect 2851 1640 2862 1674
rect 2809 1606 2862 1640
rect 1203 1512 1214 1546
rect 1248 1512 1256 1546
rect 1203 1500 1256 1512
rect 2809 1572 2817 1606
rect 2851 1572 2862 1606
rect 2809 1538 2862 1572
rect 1489 1497 1542 1509
rect 1489 1463 1497 1497
rect 1531 1463 1542 1497
rect -150 1420 -97 1432
rect -150 1386 -142 1420
rect -108 1386 -97 1420
rect -150 1352 -97 1386
rect -150 1318 -142 1352
rect -108 1318 -97 1352
rect -150 1284 -97 1318
rect -150 1250 -142 1284
rect -108 1250 -97 1284
rect -150 1232 -97 1250
rect 23 1420 79 1432
rect 23 1386 34 1420
rect 68 1386 79 1420
rect 23 1352 79 1386
rect 23 1318 34 1352
rect 68 1318 79 1352
rect 23 1284 79 1318
rect 23 1250 34 1284
rect 68 1250 79 1284
rect 23 1232 79 1250
rect 199 1420 252 1432
rect 199 1386 210 1420
rect 244 1386 252 1420
rect 199 1352 252 1386
rect 199 1318 210 1352
rect 244 1318 252 1352
rect 199 1284 252 1318
rect 199 1250 210 1284
rect 244 1250 252 1284
rect 199 1232 252 1250
rect 326 1420 379 1432
rect 326 1386 334 1420
rect 368 1386 379 1420
rect 326 1352 379 1386
rect 326 1318 334 1352
rect 368 1318 379 1352
rect 326 1284 379 1318
rect 326 1250 334 1284
rect 368 1250 379 1284
rect 326 1232 379 1250
rect 499 1420 555 1432
rect 499 1386 510 1420
rect 544 1386 555 1420
rect 499 1352 555 1386
rect 499 1318 510 1352
rect 544 1318 555 1352
rect 499 1284 555 1318
rect 499 1250 510 1284
rect 544 1250 555 1284
rect 499 1232 555 1250
rect 675 1420 731 1432
rect 675 1386 686 1420
rect 720 1386 731 1420
rect 675 1352 731 1386
rect 675 1318 686 1352
rect 720 1318 731 1352
rect 675 1284 731 1318
rect 675 1250 686 1284
rect 720 1250 731 1284
rect 675 1232 731 1250
rect 851 1420 907 1432
rect 851 1386 862 1420
rect 896 1386 907 1420
rect 851 1352 907 1386
rect 851 1318 862 1352
rect 896 1318 907 1352
rect 851 1284 907 1318
rect 851 1250 862 1284
rect 896 1250 907 1284
rect 851 1232 907 1250
rect 1027 1420 1083 1432
rect 1027 1386 1038 1420
rect 1072 1386 1083 1420
rect 1027 1352 1083 1386
rect 1027 1318 1038 1352
rect 1072 1318 1083 1352
rect 1027 1284 1083 1318
rect 1027 1250 1038 1284
rect 1072 1250 1083 1284
rect 1027 1232 1083 1250
rect 1203 1420 1256 1432
rect 1203 1386 1214 1420
rect 1248 1386 1256 1420
rect 1203 1352 1256 1386
rect 1203 1318 1214 1352
rect 1248 1318 1256 1352
rect 1203 1284 1256 1318
rect 1489 1429 1542 1463
rect 1489 1395 1497 1429
rect 1531 1395 1542 1429
rect 1489 1361 1542 1395
rect 1489 1327 1497 1361
rect 1531 1327 1542 1361
rect 1489 1309 1542 1327
rect 1662 1497 1718 1509
rect 1662 1463 1673 1497
rect 1707 1463 1718 1497
rect 1662 1429 1718 1463
rect 1662 1395 1673 1429
rect 1707 1395 1718 1429
rect 1662 1361 1718 1395
rect 1662 1327 1673 1361
rect 1707 1327 1718 1361
rect 1662 1309 1718 1327
rect 1838 1497 1894 1509
rect 1838 1463 1849 1497
rect 1883 1463 1894 1497
rect 1838 1429 1894 1463
rect 1838 1395 1849 1429
rect 1883 1395 1894 1429
rect 1838 1361 1894 1395
rect 1838 1327 1849 1361
rect 1883 1327 1894 1361
rect 1838 1309 1894 1327
rect 2014 1497 2070 1509
rect 2014 1463 2025 1497
rect 2059 1463 2070 1497
rect 2014 1429 2070 1463
rect 2014 1395 2025 1429
rect 2059 1395 2070 1429
rect 2014 1361 2070 1395
rect 2014 1327 2025 1361
rect 2059 1327 2070 1361
rect 2014 1309 2070 1327
rect 2190 1497 2246 1509
rect 2190 1463 2201 1497
rect 2235 1463 2246 1497
rect 2190 1429 2246 1463
rect 2190 1395 2201 1429
rect 2235 1395 2246 1429
rect 2190 1361 2246 1395
rect 2190 1327 2201 1361
rect 2235 1327 2246 1361
rect 2190 1309 2246 1327
rect 2366 1497 2422 1509
rect 2366 1463 2377 1497
rect 2411 1463 2422 1497
rect 2366 1429 2422 1463
rect 2366 1395 2377 1429
rect 2411 1395 2422 1429
rect 2366 1361 2422 1395
rect 2366 1327 2377 1361
rect 2411 1327 2422 1361
rect 2366 1309 2422 1327
rect 2542 1497 2595 1509
rect 2542 1463 2553 1497
rect 2587 1463 2595 1497
rect 2809 1504 2817 1538
rect 2851 1504 2862 1538
rect 2809 1492 2862 1504
rect 2982 1674 3038 1692
rect 2982 1640 2993 1674
rect 3027 1640 3038 1674
rect 2982 1606 3038 1640
rect 2982 1572 2993 1606
rect 3027 1572 3038 1606
rect 2982 1538 3038 1572
rect 2982 1504 2993 1538
rect 3027 1504 3038 1538
rect 2982 1492 3038 1504
rect 3158 1674 3214 1692
rect 3158 1640 3169 1674
rect 3203 1640 3214 1674
rect 3158 1606 3214 1640
rect 3158 1572 3169 1606
rect 3203 1572 3214 1606
rect 3158 1538 3214 1572
rect 3158 1504 3169 1538
rect 3203 1504 3214 1538
rect 3158 1492 3214 1504
rect 3334 1674 3387 1692
rect 3334 1640 3345 1674
rect 3379 1640 3387 1674
rect 3334 1606 3387 1640
rect 3334 1572 3345 1606
rect 3379 1572 3387 1606
rect 3334 1538 3387 1572
rect 3334 1504 3345 1538
rect 3379 1504 3387 1538
rect 3334 1492 3387 1504
rect 3461 1674 3514 1692
rect 3461 1640 3469 1674
rect 3503 1640 3514 1674
rect 3461 1606 3514 1640
rect 3461 1572 3469 1606
rect 3503 1572 3514 1606
rect 3461 1538 3514 1572
rect 3461 1504 3469 1538
rect 3503 1504 3514 1538
rect 3461 1492 3514 1504
rect 3634 1674 3690 1692
rect 3634 1640 3645 1674
rect 3679 1640 3690 1674
rect 3634 1606 3690 1640
rect 3634 1572 3645 1606
rect 3679 1572 3690 1606
rect 3634 1538 3690 1572
rect 3634 1504 3645 1538
rect 3679 1504 3690 1538
rect 3634 1492 3690 1504
rect 3810 1674 3866 1692
rect 3810 1640 3821 1674
rect 3855 1640 3866 1674
rect 3810 1606 3866 1640
rect 3810 1572 3821 1606
rect 3855 1572 3866 1606
rect 3810 1538 3866 1572
rect 3810 1504 3821 1538
rect 3855 1504 3866 1538
rect 3810 1492 3866 1504
rect 3986 1674 4042 1692
rect 3986 1640 3997 1674
rect 4031 1640 4042 1674
rect 3986 1606 4042 1640
rect 3986 1572 3997 1606
rect 4031 1572 4042 1606
rect 3986 1538 4042 1572
rect 3986 1504 3997 1538
rect 4031 1504 4042 1538
rect 3986 1492 4042 1504
rect 4162 1674 4215 1692
rect 4162 1640 4173 1674
rect 4207 1640 4215 1674
rect 4162 1606 4215 1640
rect 4162 1572 4173 1606
rect 4207 1572 4215 1606
rect 4162 1538 4215 1572
rect 4162 1504 4173 1538
rect 4207 1504 4215 1538
rect 4162 1492 4215 1504
rect 4289 1674 4342 1692
rect 4289 1640 4297 1674
rect 4331 1640 4342 1674
rect 4289 1606 4342 1640
rect 4289 1572 4297 1606
rect 4331 1572 4342 1606
rect 4289 1538 4342 1572
rect 4289 1504 4297 1538
rect 4331 1504 4342 1538
rect 4289 1492 4342 1504
rect 4462 1674 4518 1692
rect 4462 1640 4473 1674
rect 4507 1640 4518 1674
rect 4462 1606 4518 1640
rect 4462 1572 4473 1606
rect 4507 1572 4518 1606
rect 4462 1538 4518 1572
rect 4462 1504 4473 1538
rect 4507 1504 4518 1538
rect 4462 1492 4518 1504
rect 4638 1674 4691 1692
rect 4638 1640 4649 1674
rect 4683 1640 4691 1674
rect 4638 1606 4691 1640
rect 4638 1572 4649 1606
rect 4683 1572 4691 1606
rect 4638 1538 4691 1572
rect 4638 1504 4649 1538
rect 4683 1504 4691 1538
rect 4638 1492 4691 1504
rect 4765 1674 4818 1692
rect 4765 1640 4773 1674
rect 4807 1640 4818 1674
rect 4765 1606 4818 1640
rect 4765 1572 4773 1606
rect 4807 1572 4818 1606
rect 4765 1538 4818 1572
rect 4765 1504 4773 1538
rect 4807 1504 4818 1538
rect 4765 1492 4818 1504
rect 4938 1606 4994 1692
rect 4938 1572 4949 1606
rect 4983 1572 4994 1606
rect 4938 1538 4994 1572
rect 4938 1504 4949 1538
rect 4983 1504 4994 1538
rect 4938 1492 4994 1504
rect 5114 1674 5167 1692
rect 5114 1640 5125 1674
rect 5159 1640 5167 1674
rect 5114 1606 5167 1640
rect 5114 1572 5125 1606
rect 5159 1572 5167 1606
rect 5114 1538 5167 1572
rect 5114 1504 5125 1538
rect 5159 1504 5167 1538
rect 5114 1492 5167 1504
rect 2542 1429 2595 1463
rect 2542 1395 2553 1429
rect 2587 1395 2595 1429
rect 2542 1361 2595 1395
rect 2542 1327 2553 1361
rect 2587 1327 2595 1361
rect 2542 1309 2595 1327
rect 2809 1412 2862 1424
rect 2809 1378 2817 1412
rect 2851 1378 2862 1412
rect 2809 1344 2862 1378
rect 2809 1310 2817 1344
rect 2851 1310 2862 1344
rect 1203 1250 1214 1284
rect 1248 1250 1256 1284
rect 1203 1232 1256 1250
rect 2809 1276 2862 1310
rect 2809 1242 2817 1276
rect 2851 1242 2862 1276
rect 2809 1224 2862 1242
rect 2982 1412 3038 1424
rect 2982 1378 2993 1412
rect 3027 1378 3038 1412
rect 2982 1344 3038 1378
rect 2982 1310 2993 1344
rect 3027 1310 3038 1344
rect 2982 1276 3038 1310
rect 2982 1242 2993 1276
rect 3027 1242 3038 1276
rect 2982 1224 3038 1242
rect 3158 1412 3214 1424
rect 3158 1378 3169 1412
rect 3203 1378 3214 1412
rect 3158 1344 3214 1378
rect 3158 1310 3169 1344
rect 3203 1310 3214 1344
rect 3158 1276 3214 1310
rect 3158 1242 3169 1276
rect 3203 1242 3214 1276
rect 3158 1224 3214 1242
rect 3334 1412 3387 1424
rect 3334 1378 3345 1412
rect 3379 1378 3387 1412
rect 3334 1344 3387 1378
rect 3334 1310 3345 1344
rect 3379 1310 3387 1344
rect 3334 1276 3387 1310
rect 3334 1242 3345 1276
rect 3379 1242 3387 1276
rect 3334 1224 3387 1242
rect 3461 1412 3514 1424
rect 3461 1378 3469 1412
rect 3503 1378 3514 1412
rect 3461 1344 3514 1378
rect 3461 1310 3469 1344
rect 3503 1310 3514 1344
rect 3461 1276 3514 1310
rect 3461 1242 3469 1276
rect 3503 1242 3514 1276
rect 3461 1224 3514 1242
rect 3634 1412 3690 1424
rect 3634 1378 3645 1412
rect 3679 1378 3690 1412
rect 3634 1344 3690 1378
rect 3634 1310 3645 1344
rect 3679 1310 3690 1344
rect 3634 1276 3690 1310
rect 3634 1242 3645 1276
rect 3679 1242 3690 1276
rect 3634 1224 3690 1242
rect 3810 1412 3866 1424
rect 3810 1378 3821 1412
rect 3855 1378 3866 1412
rect 3810 1344 3866 1378
rect 3810 1310 3821 1344
rect 3855 1310 3866 1344
rect 3810 1276 3866 1310
rect 3810 1242 3821 1276
rect 3855 1242 3866 1276
rect 3810 1224 3866 1242
rect 3986 1412 4042 1424
rect 3986 1378 3997 1412
rect 4031 1378 4042 1412
rect 3986 1344 4042 1378
rect 3986 1310 3997 1344
rect 4031 1310 4042 1344
rect 3986 1276 4042 1310
rect 3986 1242 3997 1276
rect 4031 1242 4042 1276
rect 3986 1224 4042 1242
rect 4162 1412 4215 1424
rect 4162 1378 4173 1412
rect 4207 1378 4215 1412
rect 4162 1344 4215 1378
rect 4162 1310 4173 1344
rect 4207 1310 4215 1344
rect 4162 1276 4215 1310
rect 4162 1242 4173 1276
rect 4207 1242 4215 1276
rect 4162 1224 4215 1242
rect 4289 1412 4342 1424
rect 4289 1378 4297 1412
rect 4331 1378 4342 1412
rect 4289 1344 4342 1378
rect 4289 1310 4297 1344
rect 4331 1310 4342 1344
rect 4289 1276 4342 1310
rect 4289 1242 4297 1276
rect 4331 1242 4342 1276
rect 4289 1224 4342 1242
rect 4462 1412 4518 1424
rect 4462 1378 4473 1412
rect 4507 1378 4518 1412
rect 4462 1344 4518 1378
rect 4462 1310 4473 1344
rect 4507 1310 4518 1344
rect 4462 1276 4518 1310
rect 4462 1242 4473 1276
rect 4507 1242 4518 1276
rect 4462 1224 4518 1242
rect 4638 1412 4691 1424
rect 4638 1378 4649 1412
rect 4683 1378 4691 1412
rect 4638 1344 4691 1378
rect 4638 1310 4649 1344
rect 4683 1310 4691 1344
rect 4638 1276 4691 1310
rect 4638 1242 4649 1276
rect 4683 1242 4691 1276
rect 4638 1224 4691 1242
rect 4765 1412 4818 1424
rect 4765 1378 4773 1412
rect 4807 1378 4818 1412
rect 4765 1344 4818 1378
rect 4765 1310 4773 1344
rect 4807 1310 4818 1344
rect 4765 1276 4818 1310
rect 4765 1242 4773 1276
rect 4807 1242 4818 1276
rect 4765 1224 4818 1242
rect 4938 1412 4994 1424
rect 4938 1378 4949 1412
rect 4983 1378 4994 1412
rect 4938 1344 4994 1378
rect 4938 1310 4949 1344
rect 4983 1310 4994 1344
rect 4938 1276 4994 1310
rect 4938 1242 4949 1276
rect 4983 1242 4994 1276
rect 4938 1224 4994 1242
rect 5114 1412 5167 1424
rect 5114 1378 5125 1412
rect 5159 1378 5167 1412
rect 5114 1344 5167 1378
rect 5114 1310 5125 1344
rect 5159 1310 5167 1344
rect 5114 1276 5167 1310
rect 5114 1242 5125 1276
rect 5159 1242 5167 1276
rect 5114 1224 5167 1242
rect -150 1030 -97 1048
rect -150 996 -142 1030
rect -108 996 -97 1030
rect -150 962 -97 996
rect -150 928 -142 962
rect -108 928 -97 962
rect -150 894 -97 928
rect -150 860 -142 894
rect -108 860 -97 894
rect -150 848 -97 860
rect 23 1030 79 1048
rect 23 996 34 1030
rect 68 996 79 1030
rect 23 962 79 996
rect 23 928 34 962
rect 68 928 79 962
rect 23 894 79 928
rect 23 860 34 894
rect 68 860 79 894
rect 23 848 79 860
rect 199 1030 252 1048
rect 199 996 210 1030
rect 244 996 252 1030
rect 199 962 252 996
rect 199 928 210 962
rect 244 928 252 962
rect 199 894 252 928
rect 199 860 210 894
rect 244 860 252 894
rect 199 848 252 860
rect 326 1030 379 1048
rect 326 996 334 1030
rect 368 996 379 1030
rect 326 962 379 996
rect 326 928 334 962
rect 368 928 379 962
rect 326 894 379 928
rect 326 860 334 894
rect 368 860 379 894
rect 326 848 379 860
rect 499 1030 555 1048
rect 499 996 510 1030
rect 544 996 555 1030
rect 499 962 555 996
rect 499 928 510 962
rect 544 928 555 962
rect 499 894 555 928
rect 499 860 510 894
rect 544 860 555 894
rect 499 848 555 860
rect 675 1030 731 1048
rect 675 996 686 1030
rect 720 996 731 1030
rect 675 962 731 996
rect 675 928 686 962
rect 720 928 731 962
rect 675 894 731 928
rect 675 860 686 894
rect 720 860 731 894
rect 675 848 731 860
rect 851 1030 904 1048
rect 851 996 862 1030
rect 896 996 904 1030
rect 851 962 904 996
rect 851 928 862 962
rect 896 928 904 962
rect 851 894 904 928
rect 851 860 862 894
rect 896 860 904 894
rect 851 848 904 860
rect 978 1030 1031 1048
rect 978 996 986 1030
rect 1020 996 1031 1030
rect 978 962 1031 996
rect 978 928 986 962
rect 1020 928 1031 962
rect 978 894 1031 928
rect 978 860 986 894
rect 1020 860 1031 894
rect 978 848 1031 860
rect 1151 1030 1204 1048
rect 1151 996 1162 1030
rect 1196 996 1204 1030
rect 1151 962 1204 996
rect 2809 1038 2862 1056
rect 2809 1004 2817 1038
rect 2851 1004 2862 1038
rect 1151 928 1162 962
rect 1196 928 1204 962
rect 1151 894 1204 928
rect 1151 860 1162 894
rect 1196 860 1204 894
rect 1151 848 1204 860
rect 1456 956 1509 974
rect 1456 922 1464 956
rect 1498 922 1509 956
rect 1456 888 1509 922
rect 1456 854 1464 888
rect 1498 854 1509 888
rect 1456 820 1509 854
rect 1456 786 1464 820
rect 1498 786 1509 820
rect -150 768 -97 780
rect -150 734 -142 768
rect -108 734 -97 768
rect -150 700 -97 734
rect -150 666 -142 700
rect -108 666 -97 700
rect -150 632 -97 666
rect -150 598 -142 632
rect -108 598 -97 632
rect -150 580 -97 598
rect 23 768 79 780
rect 23 734 34 768
rect 68 734 79 768
rect 23 700 79 734
rect 23 666 34 700
rect 68 666 79 700
rect 23 632 79 666
rect 23 598 34 632
rect 68 598 79 632
rect 23 580 79 598
rect 199 768 252 780
rect 199 734 210 768
rect 244 734 252 768
rect 199 700 252 734
rect 199 666 210 700
rect 244 666 252 700
rect 199 632 252 666
rect 199 598 210 632
rect 244 598 252 632
rect 199 580 252 598
rect 326 768 379 780
rect 326 734 334 768
rect 368 734 379 768
rect 326 700 379 734
rect 326 666 334 700
rect 368 666 379 700
rect 326 632 379 666
rect 326 598 334 632
rect 368 598 379 632
rect 326 580 379 598
rect 499 768 555 780
rect 499 734 510 768
rect 544 734 555 768
rect 499 700 555 734
rect 499 666 510 700
rect 544 666 555 700
rect 499 632 555 666
rect 499 598 510 632
rect 544 598 555 632
rect 499 580 555 598
rect 675 768 731 780
rect 675 734 686 768
rect 720 734 731 768
rect 675 700 731 734
rect 675 666 686 700
rect 720 666 731 700
rect 675 632 731 666
rect 675 598 686 632
rect 720 598 731 632
rect 675 580 731 598
rect 851 768 904 780
rect 851 734 862 768
rect 896 734 904 768
rect 851 700 904 734
rect 851 666 862 700
rect 896 666 904 700
rect 851 632 904 666
rect 851 598 862 632
rect 896 598 904 632
rect 851 580 904 598
rect 978 768 1031 780
rect 978 734 986 768
rect 1020 734 1031 768
rect 978 700 1031 734
rect 978 666 986 700
rect 1020 666 1031 700
rect 978 632 1031 666
rect 978 598 986 632
rect 1020 598 1031 632
rect 978 580 1031 598
rect 1151 768 1204 780
rect 1456 774 1509 786
rect 1629 956 1685 974
rect 1629 922 1640 956
rect 1674 922 1685 956
rect 1629 888 1685 922
rect 1629 854 1640 888
rect 1674 854 1685 888
rect 1629 820 1685 854
rect 1629 786 1640 820
rect 1674 786 1685 820
rect 1629 774 1685 786
rect 1805 956 1861 974
rect 1805 922 1816 956
rect 1850 922 1861 956
rect 1805 888 1861 922
rect 1805 854 1816 888
rect 1850 854 1861 888
rect 1805 820 1861 854
rect 1805 786 1816 820
rect 1850 786 1861 820
rect 1805 774 1861 786
rect 1981 956 2037 974
rect 1981 922 1992 956
rect 2026 922 2037 956
rect 1981 888 2037 922
rect 1981 854 1992 888
rect 2026 854 2037 888
rect 1981 820 2037 854
rect 1981 786 1992 820
rect 2026 786 2037 820
rect 1981 774 2037 786
rect 2157 956 2213 974
rect 2157 922 2168 956
rect 2202 922 2213 956
rect 2157 888 2213 922
rect 2157 854 2168 888
rect 2202 854 2213 888
rect 2157 820 2213 854
rect 2157 786 2168 820
rect 2202 786 2213 820
rect 2157 774 2213 786
rect 2333 956 2389 974
rect 2333 922 2344 956
rect 2378 922 2389 956
rect 2333 888 2389 922
rect 2333 854 2344 888
rect 2378 854 2389 888
rect 2333 820 2389 854
rect 2333 786 2344 820
rect 2378 786 2389 820
rect 2333 774 2389 786
rect 2509 956 2562 974
rect 2509 922 2520 956
rect 2554 922 2562 956
rect 2509 888 2562 922
rect 2509 854 2520 888
rect 2554 854 2562 888
rect 2809 970 2862 1004
rect 2809 936 2817 970
rect 2851 936 2862 970
rect 2809 902 2862 936
rect 2809 868 2817 902
rect 2851 868 2862 902
rect 2809 856 2862 868
rect 2982 1038 3038 1056
rect 2982 1004 2993 1038
rect 3027 1004 3038 1038
rect 2982 970 3038 1004
rect 2982 936 2993 970
rect 3027 936 3038 970
rect 2982 902 3038 936
rect 2982 868 2993 902
rect 3027 868 3038 902
rect 2982 856 3038 868
rect 3158 1038 3214 1056
rect 3158 1004 3169 1038
rect 3203 1004 3214 1038
rect 3158 970 3214 1004
rect 3158 936 3169 970
rect 3203 936 3214 970
rect 3158 902 3214 936
rect 3158 868 3169 902
rect 3203 868 3214 902
rect 3158 856 3214 868
rect 3334 1038 3387 1056
rect 3334 1004 3345 1038
rect 3379 1004 3387 1038
rect 3334 970 3387 1004
rect 3334 936 3345 970
rect 3379 936 3387 970
rect 3334 902 3387 936
rect 3334 868 3345 902
rect 3379 868 3387 902
rect 3334 856 3387 868
rect 3461 1038 3514 1056
rect 3461 1004 3469 1038
rect 3503 1004 3514 1038
rect 3461 970 3514 1004
rect 3461 936 3469 970
rect 3503 936 3514 970
rect 3461 902 3514 936
rect 3461 868 3469 902
rect 3503 868 3514 902
rect 3461 856 3514 868
rect 3634 1038 3690 1056
rect 3634 1004 3645 1038
rect 3679 1004 3690 1038
rect 3634 970 3690 1004
rect 3634 936 3645 970
rect 3679 936 3690 970
rect 3634 902 3690 936
rect 3634 868 3645 902
rect 3679 868 3690 902
rect 3634 856 3690 868
rect 3810 1038 3863 1056
rect 3810 1004 3821 1038
rect 3855 1004 3863 1038
rect 3810 970 3863 1004
rect 3810 936 3821 970
rect 3855 936 3863 970
rect 3810 902 3863 936
rect 3810 868 3821 902
rect 3855 868 3863 902
rect 3810 856 3863 868
rect 3937 1038 3990 1056
rect 3937 1004 3945 1038
rect 3979 1004 3990 1038
rect 3937 970 3990 1004
rect 3937 936 3945 970
rect 3979 936 3990 970
rect 3937 902 3990 936
rect 3937 868 3945 902
rect 3979 868 3990 902
rect 3937 856 3990 868
rect 4110 1038 4166 1056
rect 4110 1004 4121 1038
rect 4155 1004 4166 1038
rect 4110 970 4166 1004
rect 4110 936 4121 970
rect 4155 936 4166 970
rect 4110 902 4166 936
rect 4110 868 4121 902
rect 4155 868 4166 902
rect 4110 856 4166 868
rect 4286 1038 4342 1056
rect 4286 1004 4297 1038
rect 4331 1004 4342 1038
rect 4286 970 4342 1004
rect 4286 936 4297 970
rect 4331 936 4342 970
rect 4286 902 4342 936
rect 4286 868 4297 902
rect 4331 868 4342 902
rect 4286 856 4342 868
rect 4462 1038 4518 1056
rect 4462 1004 4473 1038
rect 4507 1004 4518 1038
rect 4462 970 4518 1004
rect 4462 936 4473 970
rect 4507 936 4518 970
rect 4462 902 4518 936
rect 4462 868 4473 902
rect 4507 868 4518 902
rect 4462 856 4518 868
rect 4638 1038 4691 1056
rect 4638 1004 4649 1038
rect 4683 1004 4691 1038
rect 4638 970 4691 1004
rect 4638 936 4649 970
rect 4683 936 4691 970
rect 4638 902 4691 936
rect 4638 868 4649 902
rect 4683 868 4691 902
rect 4638 856 4691 868
rect 4765 1038 4818 1056
rect 4765 1004 4773 1038
rect 4807 1004 4818 1038
rect 4765 970 4818 1004
rect 4765 936 4773 970
rect 4807 936 4818 970
rect 4765 902 4818 936
rect 4765 868 4773 902
rect 4807 868 4818 902
rect 4765 856 4818 868
rect 4938 1038 4994 1056
rect 4938 1004 4949 1038
rect 4983 1004 4994 1038
rect 4938 970 4994 1004
rect 4938 936 4949 970
rect 4983 936 4994 970
rect 4938 902 4994 936
rect 4938 868 4949 902
rect 4983 868 4994 902
rect 4938 856 4994 868
rect 5114 1038 5167 1056
rect 5114 1004 5125 1038
rect 5159 1004 5167 1038
rect 5114 970 5167 1004
rect 5114 936 5125 970
rect 5159 936 5167 970
rect 5114 902 5167 936
rect 5114 868 5125 902
rect 5159 868 5167 902
rect 5114 856 5167 868
rect 2509 820 2562 854
rect 2509 786 2520 820
rect 2554 786 2562 820
rect 2509 774 2562 786
rect 2809 776 2862 788
rect 1151 734 1162 768
rect 1196 734 1204 768
rect 1151 700 1204 734
rect 2809 742 2817 776
rect 2851 742 2862 776
rect 2809 708 2862 742
rect 1151 666 1162 700
rect 1196 666 1204 700
rect 1151 632 1204 666
rect 1151 598 1162 632
rect 1196 598 1204 632
rect 1151 580 1204 598
rect 1456 688 1509 706
rect 1456 654 1464 688
rect 1498 654 1509 688
rect 1456 620 1509 654
rect 1456 586 1464 620
rect 1498 586 1509 620
rect 1456 552 1509 586
rect 1456 518 1464 552
rect 1498 518 1509 552
rect 1456 506 1509 518
rect 1629 688 1685 706
rect 1629 654 1640 688
rect 1674 654 1685 688
rect 1629 620 1685 654
rect 1629 586 1640 620
rect 1674 586 1685 620
rect 1629 552 1685 586
rect 1629 518 1640 552
rect 1674 518 1685 552
rect 1629 506 1685 518
rect 1805 688 1861 706
rect 1805 654 1816 688
rect 1850 654 1861 688
rect 1805 620 1861 654
rect 1805 586 1816 620
rect 1850 586 1861 620
rect 1805 552 1861 586
rect 1805 518 1816 552
rect 1850 518 1861 552
rect 1805 506 1861 518
rect 1981 688 2037 706
rect 1981 654 1992 688
rect 2026 654 2037 688
rect 1981 620 2037 654
rect 1981 586 1992 620
rect 2026 586 2037 620
rect 1981 552 2037 586
rect 1981 518 1992 552
rect 2026 518 2037 552
rect 1981 506 2037 518
rect 2157 688 2213 706
rect 2157 654 2168 688
rect 2202 654 2213 688
rect 2157 620 2213 654
rect 2157 586 2168 620
rect 2202 586 2213 620
rect 2157 552 2213 586
rect 2157 518 2168 552
rect 2202 518 2213 552
rect 2157 506 2213 518
rect 2333 688 2389 706
rect 2333 654 2344 688
rect 2378 654 2389 688
rect 2333 620 2389 654
rect 2333 586 2344 620
rect 2378 586 2389 620
rect 2333 552 2389 586
rect 2333 518 2344 552
rect 2378 518 2389 552
rect 2333 506 2389 518
rect 2509 688 2562 706
rect 2509 654 2520 688
rect 2554 654 2562 688
rect 2509 620 2562 654
rect 2509 586 2520 620
rect 2554 586 2562 620
rect 2809 674 2817 708
rect 2851 674 2862 708
rect 2809 640 2862 674
rect 2809 606 2817 640
rect 2851 606 2862 640
rect 2809 588 2862 606
rect 2982 776 3038 788
rect 2982 742 2993 776
rect 3027 742 3038 776
rect 2982 708 3038 742
rect 2982 674 2993 708
rect 3027 674 3038 708
rect 2982 640 3038 674
rect 2982 606 2993 640
rect 3027 606 3038 640
rect 2982 588 3038 606
rect 3158 776 3214 788
rect 3158 742 3169 776
rect 3203 742 3214 776
rect 3158 708 3214 742
rect 3158 674 3169 708
rect 3203 674 3214 708
rect 3158 640 3214 674
rect 3158 606 3169 640
rect 3203 606 3214 640
rect 3158 588 3214 606
rect 3334 776 3387 788
rect 3334 742 3345 776
rect 3379 742 3387 776
rect 3334 708 3387 742
rect 3334 674 3345 708
rect 3379 674 3387 708
rect 3334 640 3387 674
rect 3334 606 3345 640
rect 3379 606 3387 640
rect 3334 588 3387 606
rect 3461 776 3514 788
rect 3461 742 3469 776
rect 3503 742 3514 776
rect 3461 708 3514 742
rect 3461 674 3469 708
rect 3503 674 3514 708
rect 3461 640 3514 674
rect 3461 606 3469 640
rect 3503 606 3514 640
rect 3461 588 3514 606
rect 3634 776 3690 788
rect 3634 742 3645 776
rect 3679 742 3690 776
rect 3634 708 3690 742
rect 3634 674 3645 708
rect 3679 674 3690 708
rect 3634 640 3690 674
rect 3634 606 3645 640
rect 3679 606 3690 640
rect 3634 588 3690 606
rect 3810 776 3863 788
rect 3810 742 3821 776
rect 3855 742 3863 776
rect 3810 708 3863 742
rect 3810 674 3821 708
rect 3855 674 3863 708
rect 3810 640 3863 674
rect 3810 606 3821 640
rect 3855 606 3863 640
rect 3810 588 3863 606
rect 3937 776 3990 788
rect 3937 742 3945 776
rect 3979 742 3990 776
rect 3937 708 3990 742
rect 3937 674 3945 708
rect 3979 674 3990 708
rect 3937 640 3990 674
rect 3937 606 3945 640
rect 3979 606 3990 640
rect 3937 588 3990 606
rect 4110 776 4166 788
rect 4110 742 4121 776
rect 4155 742 4166 776
rect 4110 708 4166 742
rect 4110 674 4121 708
rect 4155 674 4166 708
rect 4110 640 4166 674
rect 4110 606 4121 640
rect 4155 606 4166 640
rect 4110 588 4166 606
rect 4286 776 4342 788
rect 4286 742 4297 776
rect 4331 742 4342 776
rect 4286 708 4342 742
rect 4286 674 4297 708
rect 4331 674 4342 708
rect 4286 640 4342 674
rect 4286 606 4297 640
rect 4331 606 4342 640
rect 4286 588 4342 606
rect 4462 776 4518 788
rect 4462 742 4473 776
rect 4507 742 4518 776
rect 4462 708 4518 742
rect 4462 674 4473 708
rect 4507 674 4518 708
rect 4462 640 4518 674
rect 4462 606 4473 640
rect 4507 606 4518 640
rect 4462 588 4518 606
rect 4638 776 4691 788
rect 4638 742 4649 776
rect 4683 742 4691 776
rect 4638 708 4691 742
rect 4638 674 4649 708
rect 4683 674 4691 708
rect 4638 640 4691 674
rect 4638 606 4649 640
rect 4683 606 4691 640
rect 4638 588 4691 606
rect 4765 776 4818 788
rect 4765 742 4773 776
rect 4807 742 4818 776
rect 4765 708 4818 742
rect 4765 674 4773 708
rect 4807 674 4818 708
rect 4765 640 4818 674
rect 4765 606 4773 640
rect 4807 606 4818 640
rect 4765 588 4818 606
rect 4938 776 4994 788
rect 4938 742 4949 776
rect 4983 742 4994 776
rect 4938 708 4994 742
rect 4938 674 4949 708
rect 4983 674 4994 708
rect 4938 640 4994 674
rect 4938 606 4949 640
rect 4983 606 4994 640
rect 4938 588 4994 606
rect 5114 776 5167 788
rect 5114 742 5125 776
rect 5159 742 5167 776
rect 5114 708 5167 742
rect 5114 674 5125 708
rect 5159 674 5167 708
rect 5114 640 5167 674
rect 5114 606 5125 640
rect 5159 606 5167 640
rect 5114 588 5167 606
rect 2509 552 2562 586
rect 2509 518 2520 552
rect 2554 518 2562 552
rect 2509 506 2562 518
<< mvndiffc >>
rect 2106 3520 2140 3554
rect 2106 3452 2140 3486
rect 2282 3520 2316 3554
rect 2282 3452 2316 3486
rect 1497 2133 1531 2167
rect 1497 2065 1531 2099
rect 1673 2133 1707 2167
rect 1673 2065 1707 2099
rect 1849 2133 1883 2167
rect 1849 2065 1883 2099
rect 2025 2133 2059 2167
rect 2025 2065 2059 2099
rect 2201 2133 2235 2167
rect 2201 2065 2235 2099
rect 2377 2133 2411 2167
rect 2377 2065 2411 2099
rect 2553 2133 2587 2167
rect 2553 2065 2587 2099
rect -142 1978 -108 2012
rect -142 1910 -108 1944
rect 34 1978 68 2012
rect 34 1910 68 1944
rect 210 1978 244 2012
rect 210 1910 244 1944
rect 334 1978 368 2012
rect 334 1910 368 1944
rect 510 1978 544 2012
rect 510 1910 544 1944
rect 686 1978 720 2012
rect 686 1910 720 1944
rect 862 1978 896 2012
rect 862 1910 896 1944
rect 1038 1978 1072 2012
rect 1038 1910 1072 1944
rect 1214 1978 1248 2012
rect 1214 1910 1248 1944
rect 2817 1970 2851 2004
rect 2817 1902 2851 1936
rect 2993 1970 3027 2004
rect 2993 1902 3027 1936
rect 3169 1970 3203 2004
rect 3169 1902 3203 1936
rect 3345 1970 3379 2004
rect 3345 1902 3379 1936
rect 3469 1970 3503 2004
rect 3469 1902 3503 1936
rect 3821 1970 3855 2004
rect 3821 1902 3855 1936
rect 4173 1970 4207 2004
rect 4173 1902 4207 1936
rect 4297 1970 4331 2004
rect 4297 1902 4331 1936
rect 4649 1970 4683 2004
rect 4649 1902 4683 1936
rect 4773 1970 4807 2004
rect 4773 1902 4807 1936
rect 4949 1970 4983 2004
rect 4949 1902 4983 1936
rect 5125 1970 5159 2004
rect 5125 1902 5159 1936
rect -142 336 -108 370
rect -142 268 -108 302
rect 210 336 244 370
rect 210 268 244 302
rect 334 336 368 370
rect 334 268 368 302
rect 510 336 544 370
rect 510 268 544 302
rect 686 336 720 370
rect 686 268 720 302
rect 862 336 896 370
rect 862 268 896 302
rect 986 336 1020 370
rect 986 268 1020 302
rect 1162 336 1196 370
rect 1162 268 1196 302
rect 2817 344 2851 378
rect 2817 276 2851 310
rect 2993 344 3027 378
rect 2993 276 3027 310
rect 3169 344 3203 378
rect 3169 276 3203 310
rect 3345 344 3379 378
rect 3345 276 3379 310
rect 3469 344 3503 378
rect 3469 276 3503 310
rect 3821 344 3855 378
rect 3821 276 3855 310
rect 3945 344 3979 378
rect 3945 276 3979 310
rect 4297 344 4331 378
rect 4297 276 4331 310
rect 4649 344 4683 378
rect 4649 276 4683 310
rect 4773 344 4807 378
rect 4773 276 4807 310
rect 5125 344 5159 378
rect 5125 276 5159 310
rect 1464 184 1498 218
rect 1464 116 1498 150
rect 1640 184 1674 218
rect 1640 116 1674 150
rect 1816 184 1850 218
rect 1816 116 1850 150
rect 1992 184 2026 218
rect 1992 116 2026 150
rect 2168 184 2202 218
rect 2168 116 2202 150
rect 2344 184 2378 218
rect 2344 116 2378 150
rect 2520 184 2554 218
rect 2520 116 2554 150
<< mvpdiffc >>
rect 2106 3190 2140 3224
rect 2106 3122 2140 3156
rect 2106 3054 2140 3088
rect 2282 3190 2316 3224
rect 2282 3122 2316 3156
rect 2282 3054 2316 3088
rect 2106 2928 2140 2962
rect 2106 2860 2140 2894
rect 2106 2792 2140 2826
rect 2282 2928 2316 2962
rect 2282 2860 2316 2894
rect 2282 2792 2316 2826
rect 1497 1731 1531 1765
rect -142 1648 -108 1682
rect -142 1580 -108 1614
rect -142 1512 -108 1546
rect 34 1580 68 1614
rect 34 1512 68 1546
rect 210 1648 244 1682
rect 210 1580 244 1614
rect 210 1512 244 1546
rect 334 1648 368 1682
rect 334 1580 368 1614
rect 334 1512 368 1546
rect 510 1648 544 1682
rect 510 1580 544 1614
rect 510 1512 544 1546
rect 686 1648 720 1682
rect 686 1580 720 1614
rect 686 1512 720 1546
rect 862 1648 896 1682
rect 862 1580 896 1614
rect 862 1512 896 1546
rect 1038 1580 1072 1614
rect 1038 1512 1072 1546
rect 1214 1648 1248 1682
rect 1214 1580 1248 1614
rect 1497 1663 1531 1697
rect 1497 1595 1531 1629
rect 1673 1731 1707 1765
rect 1673 1663 1707 1697
rect 1673 1595 1707 1629
rect 1849 1731 1883 1765
rect 1849 1663 1883 1697
rect 1849 1595 1883 1629
rect 2025 1731 2059 1765
rect 2025 1663 2059 1697
rect 2025 1595 2059 1629
rect 2201 1731 2235 1765
rect 2201 1663 2235 1697
rect 2201 1595 2235 1629
rect 2377 1731 2411 1765
rect 2377 1663 2411 1697
rect 2377 1595 2411 1629
rect 2553 1731 2587 1765
rect 2553 1663 2587 1697
rect 2553 1595 2587 1629
rect 2817 1640 2851 1674
rect 1214 1512 1248 1546
rect 2817 1572 2851 1606
rect 1497 1463 1531 1497
rect -142 1386 -108 1420
rect -142 1318 -108 1352
rect -142 1250 -108 1284
rect 34 1386 68 1420
rect 34 1318 68 1352
rect 34 1250 68 1284
rect 210 1386 244 1420
rect 210 1318 244 1352
rect 210 1250 244 1284
rect 334 1386 368 1420
rect 334 1318 368 1352
rect 334 1250 368 1284
rect 510 1386 544 1420
rect 510 1318 544 1352
rect 510 1250 544 1284
rect 686 1386 720 1420
rect 686 1318 720 1352
rect 686 1250 720 1284
rect 862 1386 896 1420
rect 862 1318 896 1352
rect 862 1250 896 1284
rect 1038 1386 1072 1420
rect 1038 1318 1072 1352
rect 1038 1250 1072 1284
rect 1214 1386 1248 1420
rect 1214 1318 1248 1352
rect 1497 1395 1531 1429
rect 1497 1327 1531 1361
rect 1673 1463 1707 1497
rect 1673 1395 1707 1429
rect 1673 1327 1707 1361
rect 1849 1463 1883 1497
rect 1849 1395 1883 1429
rect 1849 1327 1883 1361
rect 2025 1463 2059 1497
rect 2025 1395 2059 1429
rect 2025 1327 2059 1361
rect 2201 1463 2235 1497
rect 2201 1395 2235 1429
rect 2201 1327 2235 1361
rect 2377 1463 2411 1497
rect 2377 1395 2411 1429
rect 2377 1327 2411 1361
rect 2553 1463 2587 1497
rect 2817 1504 2851 1538
rect 2993 1640 3027 1674
rect 2993 1572 3027 1606
rect 2993 1504 3027 1538
rect 3169 1640 3203 1674
rect 3169 1572 3203 1606
rect 3169 1504 3203 1538
rect 3345 1640 3379 1674
rect 3345 1572 3379 1606
rect 3345 1504 3379 1538
rect 3469 1640 3503 1674
rect 3469 1572 3503 1606
rect 3469 1504 3503 1538
rect 3645 1640 3679 1674
rect 3645 1572 3679 1606
rect 3645 1504 3679 1538
rect 3821 1640 3855 1674
rect 3821 1572 3855 1606
rect 3821 1504 3855 1538
rect 3997 1640 4031 1674
rect 3997 1572 4031 1606
rect 3997 1504 4031 1538
rect 4173 1640 4207 1674
rect 4173 1572 4207 1606
rect 4173 1504 4207 1538
rect 4297 1640 4331 1674
rect 4297 1572 4331 1606
rect 4297 1504 4331 1538
rect 4473 1640 4507 1674
rect 4473 1572 4507 1606
rect 4473 1504 4507 1538
rect 4649 1640 4683 1674
rect 4649 1572 4683 1606
rect 4649 1504 4683 1538
rect 4773 1640 4807 1674
rect 4773 1572 4807 1606
rect 4773 1504 4807 1538
rect 4949 1572 4983 1606
rect 4949 1504 4983 1538
rect 5125 1640 5159 1674
rect 5125 1572 5159 1606
rect 5125 1504 5159 1538
rect 2553 1395 2587 1429
rect 2553 1327 2587 1361
rect 2817 1378 2851 1412
rect 2817 1310 2851 1344
rect 1214 1250 1248 1284
rect 2817 1242 2851 1276
rect 2993 1378 3027 1412
rect 2993 1310 3027 1344
rect 2993 1242 3027 1276
rect 3169 1378 3203 1412
rect 3169 1310 3203 1344
rect 3169 1242 3203 1276
rect 3345 1378 3379 1412
rect 3345 1310 3379 1344
rect 3345 1242 3379 1276
rect 3469 1378 3503 1412
rect 3469 1310 3503 1344
rect 3469 1242 3503 1276
rect 3645 1378 3679 1412
rect 3645 1310 3679 1344
rect 3645 1242 3679 1276
rect 3821 1378 3855 1412
rect 3821 1310 3855 1344
rect 3821 1242 3855 1276
rect 3997 1378 4031 1412
rect 3997 1310 4031 1344
rect 3997 1242 4031 1276
rect 4173 1378 4207 1412
rect 4173 1310 4207 1344
rect 4173 1242 4207 1276
rect 4297 1378 4331 1412
rect 4297 1310 4331 1344
rect 4297 1242 4331 1276
rect 4473 1378 4507 1412
rect 4473 1310 4507 1344
rect 4473 1242 4507 1276
rect 4649 1378 4683 1412
rect 4649 1310 4683 1344
rect 4649 1242 4683 1276
rect 4773 1378 4807 1412
rect 4773 1310 4807 1344
rect 4773 1242 4807 1276
rect 4949 1378 4983 1412
rect 4949 1310 4983 1344
rect 4949 1242 4983 1276
rect 5125 1378 5159 1412
rect 5125 1310 5159 1344
rect 5125 1242 5159 1276
rect -142 996 -108 1030
rect -142 928 -108 962
rect -142 860 -108 894
rect 34 996 68 1030
rect 34 928 68 962
rect 34 860 68 894
rect 210 996 244 1030
rect 210 928 244 962
rect 210 860 244 894
rect 334 996 368 1030
rect 334 928 368 962
rect 334 860 368 894
rect 510 996 544 1030
rect 510 928 544 962
rect 510 860 544 894
rect 686 996 720 1030
rect 686 928 720 962
rect 686 860 720 894
rect 862 996 896 1030
rect 862 928 896 962
rect 862 860 896 894
rect 986 996 1020 1030
rect 986 928 1020 962
rect 986 860 1020 894
rect 1162 996 1196 1030
rect 2817 1004 2851 1038
rect 1162 928 1196 962
rect 1162 860 1196 894
rect 1464 922 1498 956
rect 1464 854 1498 888
rect 1464 786 1498 820
rect -142 734 -108 768
rect -142 666 -108 700
rect -142 598 -108 632
rect 34 734 68 768
rect 34 666 68 700
rect 34 598 68 632
rect 210 734 244 768
rect 210 666 244 700
rect 210 598 244 632
rect 334 734 368 768
rect 334 666 368 700
rect 334 598 368 632
rect 510 734 544 768
rect 510 666 544 700
rect 510 598 544 632
rect 686 734 720 768
rect 686 666 720 700
rect 686 598 720 632
rect 862 734 896 768
rect 862 666 896 700
rect 862 598 896 632
rect 986 734 1020 768
rect 986 666 1020 700
rect 986 598 1020 632
rect 1640 922 1674 956
rect 1640 854 1674 888
rect 1640 786 1674 820
rect 1816 922 1850 956
rect 1816 854 1850 888
rect 1816 786 1850 820
rect 1992 922 2026 956
rect 1992 854 2026 888
rect 1992 786 2026 820
rect 2168 922 2202 956
rect 2168 854 2202 888
rect 2168 786 2202 820
rect 2344 922 2378 956
rect 2344 854 2378 888
rect 2344 786 2378 820
rect 2520 922 2554 956
rect 2520 854 2554 888
rect 2817 936 2851 970
rect 2817 868 2851 902
rect 2993 1004 3027 1038
rect 2993 936 3027 970
rect 2993 868 3027 902
rect 3169 1004 3203 1038
rect 3169 936 3203 970
rect 3169 868 3203 902
rect 3345 1004 3379 1038
rect 3345 936 3379 970
rect 3345 868 3379 902
rect 3469 1004 3503 1038
rect 3469 936 3503 970
rect 3469 868 3503 902
rect 3645 1004 3679 1038
rect 3645 936 3679 970
rect 3645 868 3679 902
rect 3821 1004 3855 1038
rect 3821 936 3855 970
rect 3821 868 3855 902
rect 3945 1004 3979 1038
rect 3945 936 3979 970
rect 3945 868 3979 902
rect 4121 1004 4155 1038
rect 4121 936 4155 970
rect 4121 868 4155 902
rect 4297 1004 4331 1038
rect 4297 936 4331 970
rect 4297 868 4331 902
rect 4473 1004 4507 1038
rect 4473 936 4507 970
rect 4473 868 4507 902
rect 4649 1004 4683 1038
rect 4649 936 4683 970
rect 4649 868 4683 902
rect 4773 1004 4807 1038
rect 4773 936 4807 970
rect 4773 868 4807 902
rect 4949 1004 4983 1038
rect 4949 936 4983 970
rect 4949 868 4983 902
rect 5125 1004 5159 1038
rect 5125 936 5159 970
rect 5125 868 5159 902
rect 2520 786 2554 820
rect 1162 734 1196 768
rect 2817 742 2851 776
rect 1162 666 1196 700
rect 1162 598 1196 632
rect 1464 654 1498 688
rect 1464 586 1498 620
rect 1464 518 1498 552
rect 1640 654 1674 688
rect 1640 586 1674 620
rect 1640 518 1674 552
rect 1816 654 1850 688
rect 1816 586 1850 620
rect 1816 518 1850 552
rect 1992 654 2026 688
rect 1992 586 2026 620
rect 1992 518 2026 552
rect 2168 654 2202 688
rect 2168 586 2202 620
rect 2168 518 2202 552
rect 2344 654 2378 688
rect 2344 586 2378 620
rect 2344 518 2378 552
rect 2520 654 2554 688
rect 2520 586 2554 620
rect 2817 674 2851 708
rect 2817 606 2851 640
rect 2993 742 3027 776
rect 2993 674 3027 708
rect 2993 606 3027 640
rect 3169 742 3203 776
rect 3169 674 3203 708
rect 3169 606 3203 640
rect 3345 742 3379 776
rect 3345 674 3379 708
rect 3345 606 3379 640
rect 3469 742 3503 776
rect 3469 674 3503 708
rect 3469 606 3503 640
rect 3645 742 3679 776
rect 3645 674 3679 708
rect 3645 606 3679 640
rect 3821 742 3855 776
rect 3821 674 3855 708
rect 3821 606 3855 640
rect 3945 742 3979 776
rect 3945 674 3979 708
rect 3945 606 3979 640
rect 4121 742 4155 776
rect 4121 674 4155 708
rect 4121 606 4155 640
rect 4297 742 4331 776
rect 4297 674 4331 708
rect 4297 606 4331 640
rect 4473 742 4507 776
rect 4473 674 4507 708
rect 4473 606 4507 640
rect 4649 742 4683 776
rect 4649 674 4683 708
rect 4649 606 4683 640
rect 4773 742 4807 776
rect 4773 674 4807 708
rect 4773 606 4807 640
rect 4949 742 4983 776
rect 4949 674 4983 708
rect 4949 606 4983 640
rect 5125 742 5159 776
rect 5125 674 5159 708
rect 5125 606 5159 640
rect 2520 518 2554 552
<< mvpsubdiff >>
rect 2095 3677 2119 3711
rect 2153 3677 2253 3711
rect 2287 3677 2311 3711
rect 2784 2251 2840 2285
rect 2874 2251 2908 2285
rect 2942 2251 2976 2285
rect 3010 2251 3044 2285
rect 3078 2251 3112 2285
rect 3146 2251 3180 2285
rect 3214 2251 3248 2285
rect 3282 2251 3316 2285
rect 3350 2251 3384 2285
rect 3418 2251 3452 2285
rect 3486 2251 3520 2285
rect 3554 2251 3588 2285
rect 3622 2251 3656 2285
rect 3690 2251 3714 2285
rect 2784 2211 3714 2251
rect 306 2112 371 2146
rect 405 2112 439 2146
rect 473 2112 507 2146
rect 541 2112 575 2146
rect 609 2112 643 2146
rect 677 2112 711 2146
rect 745 2112 779 2146
rect 813 2112 847 2146
rect 881 2112 915 2146
rect 949 2112 983 2146
rect 1017 2112 1051 2146
rect 1085 2112 1119 2146
rect 1153 2112 1187 2146
rect 1221 2112 1255 2146
rect 1289 2112 1313 2146
rect 2784 2177 2840 2211
rect 2874 2177 2908 2211
rect 2942 2177 2976 2211
rect 3010 2177 3044 2211
rect 3078 2177 3112 2211
rect 3146 2177 3180 2211
rect 3214 2177 3248 2211
rect 3282 2177 3316 2211
rect 3350 2177 3384 2211
rect 3418 2177 3452 2211
rect 3486 2177 3520 2211
rect 3554 2177 3588 2211
rect 3622 2177 3656 2211
rect 3690 2177 3714 2211
rect 2784 2138 3714 2177
rect 2784 2104 2868 2138
rect 2902 2104 2936 2138
rect 2970 2104 3004 2138
rect 3038 2104 3072 2138
rect 3106 2104 3140 2138
rect 3174 2104 3208 2138
rect 3242 2104 3276 2138
rect 3310 2104 3344 2138
rect 3378 2104 3412 2138
rect 3446 2104 3480 2138
rect 3514 2104 3548 2138
rect 3582 2104 3616 2138
rect 3650 2104 3684 2138
rect 3718 2104 3752 2138
rect 3786 2104 3820 2138
rect 3854 2104 3888 2138
rect 3922 2104 3956 2138
rect 3990 2104 4024 2138
rect 4058 2104 4092 2138
rect 4126 2104 4160 2138
rect 4194 2104 4228 2138
rect 4262 2104 4296 2138
rect 4330 2104 4364 2138
rect 4398 2104 4432 2138
rect 4466 2104 4500 2138
rect 4534 2104 4568 2138
rect 4602 2104 4636 2138
rect 4670 2104 4704 2138
rect 4738 2104 4772 2138
rect 4806 2104 4840 2138
rect 4874 2104 4908 2138
rect 4942 2104 4976 2138
rect 5010 2104 5044 2138
rect 5078 2104 5112 2138
rect 5146 2104 5170 2138
rect 317 117 373 151
rect 407 117 441 151
rect 475 117 509 151
rect 543 117 577 151
rect 611 117 645 151
rect 679 117 713 151
rect 747 117 781 151
rect 815 117 849 151
rect 883 117 917 151
rect 951 117 985 151
rect 1019 117 1053 151
rect 1087 117 1121 151
rect 1155 117 1189 151
rect 1223 117 1247 151
rect 2805 142 2865 176
rect 2899 142 2933 176
rect 2967 142 3001 176
rect 3035 142 3069 176
rect 3103 142 3137 176
rect 3171 142 3205 176
rect 3239 142 3273 176
rect 3307 142 3341 176
rect 3375 142 3409 176
rect 3443 142 3477 176
rect 3511 142 3545 176
rect 3579 142 3613 176
rect 3647 142 3681 176
rect 3715 142 3749 176
rect 3783 142 3817 176
rect 3851 142 3885 176
rect 3919 142 3953 176
rect 3987 142 4021 176
rect 4055 142 4089 176
rect 4123 142 4157 176
rect 4191 142 4225 176
rect 4259 142 4293 176
rect 4327 142 4361 176
rect 4395 142 4429 176
rect 4463 142 4497 176
rect 4531 142 4565 176
rect 4599 142 4633 176
rect 4667 142 4701 176
rect 4735 142 4769 176
rect 4803 142 4837 176
rect 4871 142 4905 176
rect 4939 142 4973 176
rect 5007 142 5041 176
rect 5075 142 5109 176
rect 5143 142 5167 176
<< mvnsubdiff >>
rect 2075 2621 2099 2655
rect 2133 2621 2183 2655
rect 2217 2621 2266 2655
rect 2300 2621 2324 2655
rect 2075 2587 2324 2621
rect 2075 2553 2099 2587
rect 2133 2553 2183 2587
rect 2217 2553 2266 2587
rect 2300 2553 2324 2587
rect 353 1123 425 1157
rect 459 1123 493 1157
rect 527 1123 561 1157
rect 595 1123 629 1157
rect 663 1123 697 1157
rect 731 1123 765 1157
rect 799 1123 833 1157
rect 867 1123 901 1157
rect 935 1123 969 1157
rect 1003 1123 1037 1157
rect 1071 1123 1105 1157
rect 1139 1123 1173 1157
rect 1207 1123 1241 1157
rect 1275 1123 1309 1157
rect 1343 1123 1377 1157
rect 1411 1123 1515 1157
rect 1549 1123 1583 1157
rect 1617 1123 1651 1157
rect 1685 1123 1719 1157
rect 1753 1123 1787 1157
rect 1821 1123 1855 1157
rect 1889 1123 1923 1157
rect 1957 1123 1991 1157
rect 2025 1123 2059 1157
rect 2093 1123 2127 1157
rect 2161 1123 2195 1157
rect 2229 1123 2263 1157
rect 2297 1123 2331 1157
rect 2365 1123 2399 1157
rect 2433 1123 2467 1157
rect 2501 1123 2532 1157
rect 2809 1123 2865 1157
rect 2899 1123 2933 1157
rect 2967 1123 3001 1157
rect 3035 1123 3069 1157
rect 3103 1123 3137 1157
rect 3171 1123 3205 1157
rect 3239 1123 3273 1157
rect 3307 1123 3341 1157
rect 3375 1123 3409 1157
rect 3443 1123 3477 1157
rect 3511 1123 3545 1157
rect 3579 1123 3613 1157
rect 3647 1123 3681 1157
rect 3715 1123 3749 1157
rect 3783 1123 3817 1157
rect 3851 1123 3885 1157
rect 3919 1123 3953 1157
rect 3987 1123 4021 1157
rect 4055 1123 4089 1157
rect 4123 1123 4157 1157
rect 4191 1123 4225 1157
rect 4259 1123 4293 1157
rect 4327 1123 4361 1157
rect 4395 1123 4429 1157
rect 4463 1123 4497 1157
rect 4531 1123 4565 1157
rect 4599 1123 4633 1157
rect 4667 1123 4701 1157
rect 4735 1123 4769 1157
rect 4803 1123 4837 1157
rect 4871 1123 4905 1157
rect 4939 1123 4973 1157
rect 5007 1123 5041 1157
rect 5075 1123 5109 1157
rect 5143 1123 5167 1157
<< mvpsubdiffcont >>
rect 2119 3677 2153 3711
rect 2253 3677 2287 3711
rect 2840 2251 2874 2285
rect 2908 2251 2942 2285
rect 2976 2251 3010 2285
rect 3044 2251 3078 2285
rect 3112 2251 3146 2285
rect 3180 2251 3214 2285
rect 3248 2251 3282 2285
rect 3316 2251 3350 2285
rect 3384 2251 3418 2285
rect 3452 2251 3486 2285
rect 3520 2251 3554 2285
rect 3588 2251 3622 2285
rect 3656 2251 3690 2285
rect 371 2112 405 2146
rect 439 2112 473 2146
rect 507 2112 541 2146
rect 575 2112 609 2146
rect 643 2112 677 2146
rect 711 2112 745 2146
rect 779 2112 813 2146
rect 847 2112 881 2146
rect 915 2112 949 2146
rect 983 2112 1017 2146
rect 1051 2112 1085 2146
rect 1119 2112 1153 2146
rect 1187 2112 1221 2146
rect 1255 2112 1289 2146
rect 2840 2177 2874 2211
rect 2908 2177 2942 2211
rect 2976 2177 3010 2211
rect 3044 2177 3078 2211
rect 3112 2177 3146 2211
rect 3180 2177 3214 2211
rect 3248 2177 3282 2211
rect 3316 2177 3350 2211
rect 3384 2177 3418 2211
rect 3452 2177 3486 2211
rect 3520 2177 3554 2211
rect 3588 2177 3622 2211
rect 3656 2177 3690 2211
rect 2868 2104 2902 2138
rect 2936 2104 2970 2138
rect 3004 2104 3038 2138
rect 3072 2104 3106 2138
rect 3140 2104 3174 2138
rect 3208 2104 3242 2138
rect 3276 2104 3310 2138
rect 3344 2104 3378 2138
rect 3412 2104 3446 2138
rect 3480 2104 3514 2138
rect 3548 2104 3582 2138
rect 3616 2104 3650 2138
rect 3684 2104 3718 2138
rect 3752 2104 3786 2138
rect 3820 2104 3854 2138
rect 3888 2104 3922 2138
rect 3956 2104 3990 2138
rect 4024 2104 4058 2138
rect 4092 2104 4126 2138
rect 4160 2104 4194 2138
rect 4228 2104 4262 2138
rect 4296 2104 4330 2138
rect 4364 2104 4398 2138
rect 4432 2104 4466 2138
rect 4500 2104 4534 2138
rect 4568 2104 4602 2138
rect 4636 2104 4670 2138
rect 4704 2104 4738 2138
rect 4772 2104 4806 2138
rect 4840 2104 4874 2138
rect 4908 2104 4942 2138
rect 4976 2104 5010 2138
rect 5044 2104 5078 2138
rect 5112 2104 5146 2138
rect 373 117 407 151
rect 441 117 475 151
rect 509 117 543 151
rect 577 117 611 151
rect 645 117 679 151
rect 713 117 747 151
rect 781 117 815 151
rect 849 117 883 151
rect 917 117 951 151
rect 985 117 1019 151
rect 1053 117 1087 151
rect 1121 117 1155 151
rect 1189 117 1223 151
rect 2865 142 2899 176
rect 2933 142 2967 176
rect 3001 142 3035 176
rect 3069 142 3103 176
rect 3137 142 3171 176
rect 3205 142 3239 176
rect 3273 142 3307 176
rect 3341 142 3375 176
rect 3409 142 3443 176
rect 3477 142 3511 176
rect 3545 142 3579 176
rect 3613 142 3647 176
rect 3681 142 3715 176
rect 3749 142 3783 176
rect 3817 142 3851 176
rect 3885 142 3919 176
rect 3953 142 3987 176
rect 4021 142 4055 176
rect 4089 142 4123 176
rect 4157 142 4191 176
rect 4225 142 4259 176
rect 4293 142 4327 176
rect 4361 142 4395 176
rect 4429 142 4463 176
rect 4497 142 4531 176
rect 4565 142 4599 176
rect 4633 142 4667 176
rect 4701 142 4735 176
rect 4769 142 4803 176
rect 4837 142 4871 176
rect 4905 142 4939 176
rect 4973 142 5007 176
rect 5041 142 5075 176
rect 5109 142 5143 176
<< mvnsubdiffcont >>
rect 2099 2621 2133 2655
rect 2183 2621 2217 2655
rect 2266 2621 2300 2655
rect 2099 2553 2133 2587
rect 2183 2553 2217 2587
rect 2266 2553 2300 2587
rect 425 1123 459 1157
rect 493 1123 527 1157
rect 561 1123 595 1157
rect 629 1123 663 1157
rect 697 1123 731 1157
rect 765 1123 799 1157
rect 833 1123 867 1157
rect 901 1123 935 1157
rect 969 1123 1003 1157
rect 1037 1123 1071 1157
rect 1105 1123 1139 1157
rect 1173 1123 1207 1157
rect 1241 1123 1275 1157
rect 1309 1123 1343 1157
rect 1377 1123 1411 1157
rect 1515 1123 1549 1157
rect 1583 1123 1617 1157
rect 1651 1123 1685 1157
rect 1719 1123 1753 1157
rect 1787 1123 1821 1157
rect 1855 1123 1889 1157
rect 1923 1123 1957 1157
rect 1991 1123 2025 1157
rect 2059 1123 2093 1157
rect 2127 1123 2161 1157
rect 2195 1123 2229 1157
rect 2263 1123 2297 1157
rect 2331 1123 2365 1157
rect 2399 1123 2433 1157
rect 2467 1123 2501 1157
rect 2865 1123 2899 1157
rect 2933 1123 2967 1157
rect 3001 1123 3035 1157
rect 3069 1123 3103 1157
rect 3137 1123 3171 1157
rect 3205 1123 3239 1157
rect 3273 1123 3307 1157
rect 3341 1123 3375 1157
rect 3409 1123 3443 1157
rect 3477 1123 3511 1157
rect 3545 1123 3579 1157
rect 3613 1123 3647 1157
rect 3681 1123 3715 1157
rect 3749 1123 3783 1157
rect 3817 1123 3851 1157
rect 3885 1123 3919 1157
rect 3953 1123 3987 1157
rect 4021 1123 4055 1157
rect 4089 1123 4123 1157
rect 4157 1123 4191 1157
rect 4225 1123 4259 1157
rect 4293 1123 4327 1157
rect 4361 1123 4395 1157
rect 4429 1123 4463 1157
rect 4497 1123 4531 1157
rect 4565 1123 4599 1157
rect 4633 1123 4667 1157
rect 4701 1123 4735 1157
rect 4769 1123 4803 1157
rect 4837 1123 4871 1157
rect 4905 1123 4939 1157
rect 4973 1123 5007 1157
rect 5041 1123 5075 1157
rect 5109 1123 5143 1157
<< poly >>
rect 2151 3580 2271 3606
rect 2151 3392 2271 3440
rect 2151 3358 2195 3392
rect 2229 3358 2271 3392
rect 2151 3324 2271 3358
rect 2151 3290 2195 3324
rect 2229 3290 2271 3324
rect 2151 3242 2271 3290
rect 2151 2974 2271 3042
rect 2151 2748 2271 2774
rect 1536 2255 1670 2271
rect 1536 2221 1552 2255
rect 1586 2221 1620 2255
rect 1654 2221 1670 2255
rect 1536 2205 1670 2221
rect 2064 2255 2198 2271
rect 2064 2221 2080 2255
rect 2114 2221 2148 2255
rect 2182 2221 2198 2255
rect 2064 2205 2198 2221
rect 2246 2255 2542 2271
rect 2246 2221 2262 2255
rect 2296 2221 2338 2255
rect 2372 2221 2415 2255
rect 2449 2221 2492 2255
rect 2526 2221 2542 2255
rect 2246 2205 2542 2221
rect 1542 2179 1662 2205
rect 1718 2179 1838 2205
rect 1894 2179 2014 2205
rect 2070 2179 2190 2205
rect 2246 2179 2366 2205
rect 2422 2179 2542 2205
rect -97 2038 23 2064
rect 79 2038 199 2064
rect 379 2038 499 2064
rect 555 2038 675 2064
rect 731 2038 851 2064
rect 907 2038 1027 2064
rect 1083 2038 1203 2064
rect -97 1850 23 1898
rect -97 1816 -54 1850
rect -20 1816 23 1850
rect -97 1782 23 1816
rect -97 1748 -54 1782
rect -20 1748 23 1782
rect -97 1700 23 1748
rect 79 1850 199 1898
rect 79 1816 124 1850
rect 158 1816 199 1850
rect 79 1782 199 1816
rect 79 1748 124 1782
rect 158 1748 199 1782
rect 79 1700 199 1748
rect 379 1850 499 1898
rect 379 1816 421 1850
rect 455 1816 499 1850
rect 379 1782 499 1816
rect 379 1748 421 1782
rect 455 1748 499 1782
rect 379 1700 499 1748
rect 555 1872 675 1898
rect 731 1872 851 1898
rect 555 1850 851 1872
rect 555 1816 592 1850
rect 626 1816 779 1850
rect 813 1816 851 1850
rect 555 1782 851 1816
rect 555 1748 592 1782
rect 626 1748 779 1782
rect 813 1748 851 1782
rect 555 1726 851 1748
rect 555 1700 675 1726
rect 731 1700 851 1726
rect 907 1850 1027 1898
rect 907 1816 950 1850
rect 984 1816 1027 1850
rect 907 1782 1027 1816
rect 907 1748 950 1782
rect 984 1748 1027 1782
rect 907 1700 1027 1748
rect 1083 1850 1203 1898
rect 1083 1816 1128 1850
rect 1162 1816 1203 1850
rect 1083 1782 1203 1816
rect 1083 1748 1128 1782
rect 1162 1748 1203 1782
rect 1542 1777 1662 2039
rect 1718 1890 1838 2039
rect 1894 1971 2014 2039
rect 2070 2013 2190 2039
rect 1894 1937 2190 1971
rect 1894 1932 2114 1937
rect 2070 1903 2114 1932
rect 2148 1903 2190 1937
rect 1718 1851 2014 1890
rect 1718 1777 1838 1809
rect 1894 1777 2014 1851
rect 2070 1869 2190 1903
rect 2070 1835 2114 1869
rect 2148 1835 2190 1869
rect 2070 1777 2190 1835
rect 2246 1777 2366 2039
rect 2422 1777 2542 2039
rect 2862 2030 2982 2056
rect 3038 2030 3158 2056
rect 3214 2030 3334 2056
rect 3514 2030 3634 2056
rect 3690 2030 3810 2056
rect 3866 2030 3986 2056
rect 4042 2030 4162 2056
rect 4342 2030 4462 2056
rect 4518 2030 4638 2056
rect 4818 2030 4938 2056
rect 4994 2030 5114 2056
rect 2862 1864 2982 1890
rect 3038 1864 3158 1890
rect 2862 1842 3158 1864
rect 2862 1808 2900 1842
rect 2934 1808 3087 1842
rect 3121 1808 3158 1842
rect 1083 1700 1203 1748
rect 2862 1774 3158 1808
rect 2862 1740 2900 1774
rect 2934 1740 3087 1774
rect 3121 1740 3158 1774
rect 2862 1718 3158 1740
rect 2862 1692 2982 1718
rect 3038 1692 3158 1718
rect 3214 1842 3334 1890
rect 3214 1808 3258 1842
rect 3292 1808 3334 1842
rect 3214 1774 3334 1808
rect 3214 1740 3258 1774
rect 3292 1740 3334 1774
rect 3214 1692 3334 1740
rect 3514 1842 3634 1890
rect 3514 1808 3559 1842
rect 3593 1808 3634 1842
rect 3514 1774 3634 1808
rect 3514 1740 3559 1774
rect 3593 1740 3634 1774
rect 3514 1692 3634 1740
rect 3690 1842 3810 1890
rect 3690 1808 3730 1842
rect 3764 1808 3810 1842
rect 3690 1774 3810 1808
rect 3690 1740 3730 1774
rect 3764 1740 3810 1774
rect 3690 1692 3810 1740
rect 3866 1842 3986 1890
rect 3866 1808 3912 1842
rect 3946 1808 3986 1842
rect 3866 1774 3986 1808
rect 3866 1740 3912 1774
rect 3946 1740 3986 1774
rect 3866 1692 3986 1740
rect 4042 1842 4162 1890
rect 4042 1808 4083 1842
rect 4117 1808 4162 1842
rect 4042 1774 4162 1808
rect 4042 1740 4083 1774
rect 4117 1740 4162 1774
rect 4042 1692 4162 1740
rect 4342 1842 4462 1890
rect 4342 1808 4387 1842
rect 4421 1808 4462 1842
rect 4342 1774 4462 1808
rect 4342 1740 4387 1774
rect 4421 1740 4462 1774
rect 4342 1692 4462 1740
rect 4518 1842 4638 1890
rect 4518 1808 4558 1842
rect 4592 1808 4638 1842
rect 4518 1774 4638 1808
rect 4518 1740 4558 1774
rect 4592 1740 4638 1774
rect 4518 1692 4638 1740
rect 4818 1842 4938 1890
rect 4818 1808 4861 1842
rect 4895 1808 4938 1842
rect 4818 1774 4938 1808
rect 4818 1740 4861 1774
rect 4895 1740 4938 1774
rect 4818 1692 4938 1740
rect 4994 1842 5114 1890
rect 4994 1808 5039 1842
rect 5073 1808 5114 1842
rect 4994 1774 5114 1808
rect 4994 1740 5039 1774
rect 5073 1740 5114 1774
rect 4994 1692 5114 1740
rect 1542 1509 1662 1577
rect 1718 1509 1838 1577
rect 1894 1509 2014 1577
rect 2070 1509 2190 1577
rect 2246 1509 2366 1577
rect 2422 1509 2542 1577
rect -97 1432 23 1500
rect 79 1432 199 1500
rect 379 1432 499 1500
rect 555 1432 675 1500
rect 731 1432 851 1500
rect 907 1432 1027 1500
rect 1083 1432 1203 1500
rect 2862 1424 2982 1492
rect 3038 1424 3158 1492
rect 3214 1424 3334 1492
rect 3514 1424 3634 1492
rect 3690 1424 3810 1492
rect 3866 1424 3986 1492
rect 4042 1424 4162 1492
rect 4342 1424 4462 1492
rect 4518 1424 4638 1492
rect 4818 1424 4938 1492
rect 4994 1424 5114 1492
rect 1542 1277 1662 1309
rect 1718 1277 1838 1309
rect 1894 1277 2014 1309
rect 2070 1277 2190 1309
rect 2246 1277 2366 1309
rect 2422 1277 2542 1309
rect 1542 1261 1838 1277
rect -97 1206 23 1232
rect 79 1206 199 1232
rect 379 1206 499 1232
rect 555 1206 675 1232
rect 731 1206 851 1232
rect 907 1206 1027 1232
rect 1083 1206 1203 1232
rect 1542 1227 1558 1261
rect 1592 1227 1634 1261
rect 1668 1227 1711 1261
rect 1745 1227 1788 1261
rect 1822 1227 1838 1261
rect 1542 1211 1838 1227
rect 1888 1261 2022 1277
rect 1888 1227 1904 1261
rect 1938 1227 1972 1261
rect 2006 1227 2022 1261
rect 1888 1211 2022 1227
rect 2246 1261 2542 1277
rect 2246 1227 2262 1261
rect 2296 1227 2338 1261
rect 2372 1227 2415 1261
rect 2449 1227 2492 1261
rect 2526 1227 2542 1261
rect 2246 1211 2542 1227
rect 2862 1198 2982 1224
rect 3038 1198 3158 1224
rect 3214 1198 3334 1224
rect 3514 1198 3634 1224
rect 3690 1198 3810 1224
rect 3866 1198 3986 1224
rect 4042 1198 4162 1224
rect 4342 1198 4462 1224
rect 4518 1198 4638 1224
rect 4818 1198 4938 1224
rect 4994 1198 5114 1224
rect -97 1048 23 1074
rect 79 1048 199 1074
rect 379 1048 499 1074
rect 555 1048 675 1074
rect 731 1048 851 1074
rect 1031 1048 1151 1074
rect 1509 1056 1805 1072
rect 1509 1022 1525 1056
rect 1559 1022 1601 1056
rect 1635 1022 1678 1056
rect 1712 1022 1755 1056
rect 1789 1022 1805 1056
rect 1509 1006 1805 1022
rect 1855 1056 1989 1072
rect 1855 1022 1871 1056
rect 1905 1022 1939 1056
rect 1973 1022 1989 1056
rect 1855 1006 1989 1022
rect 2213 1056 2509 1072
rect 2862 1056 2982 1082
rect 3038 1056 3158 1082
rect 3214 1056 3334 1082
rect 3514 1056 3634 1082
rect 3690 1056 3810 1082
rect 3990 1056 4110 1082
rect 4166 1056 4286 1082
rect 4342 1056 4462 1082
rect 4518 1056 4638 1082
rect 4818 1056 4938 1082
rect 4994 1056 5114 1082
rect 2213 1022 2229 1056
rect 2263 1022 2305 1056
rect 2339 1022 2382 1056
rect 2416 1022 2459 1056
rect 2493 1022 2509 1056
rect 2213 1006 2509 1022
rect 1509 974 1629 1006
rect 1685 974 1805 1006
rect 1861 974 1981 1006
rect 2037 974 2157 1006
rect 2213 974 2333 1006
rect 2389 974 2509 1006
rect -97 780 23 848
rect 79 780 199 848
rect 379 780 499 848
rect 555 780 675 848
rect 731 780 851 848
rect 1031 780 1151 848
rect 2862 788 2982 856
rect 3038 788 3158 856
rect 3214 788 3334 856
rect 3514 788 3634 856
rect 3690 788 3810 856
rect 3990 788 4110 856
rect 4166 788 4286 856
rect 4342 788 4462 856
rect 4518 788 4638 856
rect 4818 788 4938 856
rect 4994 788 5114 856
rect 1509 706 1629 774
rect 1685 706 1805 774
rect 1861 706 1981 774
rect 2037 706 2157 774
rect 2213 706 2333 774
rect 2389 706 2509 774
rect -97 532 23 580
rect -97 498 -52 532
rect -18 498 23 532
rect -97 464 23 498
rect -97 430 -52 464
rect -18 430 23 464
rect -97 382 23 430
rect 79 532 199 580
rect 79 498 119 532
rect 153 498 199 532
rect 79 464 199 498
rect 79 430 119 464
rect 153 430 199 464
rect 79 382 199 430
rect 379 532 499 580
rect 379 498 421 532
rect 455 498 499 532
rect 379 464 499 498
rect 379 430 421 464
rect 455 430 499 464
rect 379 382 499 430
rect 555 554 675 580
rect 731 554 851 580
rect 555 532 851 554
rect 555 498 592 532
rect 626 498 779 532
rect 813 498 851 532
rect 555 464 851 498
rect 555 430 592 464
rect 626 430 779 464
rect 813 430 851 464
rect 555 408 851 430
rect 555 382 675 408
rect 731 382 851 408
rect 1031 532 1151 580
rect 1031 498 1073 532
rect 1107 498 1151 532
rect 2862 562 2982 588
rect 3038 562 3158 588
rect 2862 540 3158 562
rect 2862 506 2899 540
rect 2933 506 3086 540
rect 3120 506 3158 540
rect 1031 464 1151 498
rect 1031 430 1073 464
rect 1107 430 1151 464
rect 1031 382 1151 430
rect 1509 244 1629 506
rect 1685 474 1805 506
rect 1861 432 1981 506
rect 1685 393 1981 432
rect 2037 448 2157 506
rect 2037 414 2081 448
rect 2115 414 2157 448
rect 1685 244 1805 393
rect 2037 380 2157 414
rect 2037 351 2081 380
rect 1861 346 2081 351
rect 2115 346 2157 380
rect 1861 312 2157 346
rect 1861 244 1981 312
rect 2037 244 2157 270
rect 2213 244 2333 506
rect 2389 244 2509 506
rect 2862 472 3158 506
rect 2862 438 2899 472
rect 2933 438 3086 472
rect 3120 438 3158 472
rect 2862 416 3158 438
rect 2862 390 2982 416
rect 3038 390 3158 416
rect 3214 540 3334 588
rect 3214 506 3258 540
rect 3292 506 3334 540
rect 3214 472 3334 506
rect 3214 438 3258 472
rect 3292 438 3334 472
rect 3214 390 3334 438
rect 3514 540 3634 588
rect 3514 506 3560 540
rect 3594 506 3634 540
rect 3514 472 3634 506
rect 3514 438 3560 472
rect 3594 438 3634 472
rect 3514 390 3634 438
rect 3690 540 3810 588
rect 3690 506 3731 540
rect 3765 506 3810 540
rect 3690 472 3810 506
rect 3690 438 3731 472
rect 3765 438 3810 472
rect 3690 390 3810 438
rect 3990 540 4110 588
rect 3990 506 4035 540
rect 4069 506 4110 540
rect 3990 472 4110 506
rect 3990 438 4035 472
rect 4069 438 4110 472
rect 3990 390 4110 438
rect 4166 540 4286 588
rect 4166 506 4206 540
rect 4240 506 4286 540
rect 4166 472 4286 506
rect 4166 438 4206 472
rect 4240 438 4286 472
rect 4166 390 4286 438
rect 4342 540 4462 588
rect 4342 506 4388 540
rect 4422 506 4462 540
rect 4342 472 4462 506
rect 4342 438 4388 472
rect 4422 438 4462 472
rect 4342 390 4462 438
rect 4518 540 4638 588
rect 4518 506 4559 540
rect 4593 506 4638 540
rect 4518 472 4638 506
rect 4518 438 4559 472
rect 4593 438 4638 472
rect 4518 390 4638 438
rect 4818 540 4938 588
rect 4818 506 4864 540
rect 4898 506 4938 540
rect 4818 472 4938 506
rect 4818 438 4864 472
rect 4898 438 4938 472
rect 4818 390 4938 438
rect 4994 540 5114 588
rect 4994 506 5035 540
rect 5069 506 5114 540
rect 4994 472 5114 506
rect 4994 438 5035 472
rect 5069 438 5114 472
rect 4994 390 5114 438
rect -97 216 23 242
rect 79 216 199 242
rect 379 216 499 242
rect 555 216 675 242
rect 731 216 851 242
rect 1031 216 1151 242
rect 2862 224 2982 250
rect 3038 224 3158 250
rect 3214 224 3334 250
rect 3514 224 3634 250
rect 3690 224 3810 250
rect 3990 224 4110 250
rect 4166 224 4286 250
rect 4342 224 4462 250
rect 4518 224 4638 250
rect 4818 224 4938 250
rect 4994 224 5114 250
rect 1509 78 1629 104
rect 1685 78 1805 104
rect 1861 78 1981 104
rect 2037 78 2157 104
rect 2213 78 2333 104
rect 2389 78 2509 104
rect 1503 62 1637 78
rect 1503 28 1519 62
rect 1553 28 1587 62
rect 1621 28 1637 62
rect 1503 12 1637 28
rect 2031 62 2165 78
rect 2031 28 2047 62
rect 2081 28 2115 62
rect 2149 28 2165 62
rect 2031 12 2165 28
rect 2213 62 2509 78
rect 2213 28 2229 62
rect 2263 28 2305 62
rect 2339 28 2382 62
rect 2416 28 2459 62
rect 2493 28 2509 62
rect 2213 12 2509 28
<< polycont >>
rect 2195 3358 2229 3392
rect 2195 3290 2229 3324
rect 1552 2221 1586 2255
rect 1620 2221 1654 2255
rect 2080 2221 2114 2255
rect 2148 2221 2182 2255
rect 2262 2221 2296 2255
rect 2338 2221 2372 2255
rect 2415 2221 2449 2255
rect 2492 2221 2526 2255
rect -54 1816 -20 1850
rect -54 1748 -20 1782
rect 124 1816 158 1850
rect 124 1748 158 1782
rect 421 1816 455 1850
rect 421 1748 455 1782
rect 592 1816 626 1850
rect 779 1816 813 1850
rect 592 1748 626 1782
rect 779 1748 813 1782
rect 950 1816 984 1850
rect 950 1748 984 1782
rect 1128 1816 1162 1850
rect 1128 1748 1162 1782
rect 2114 1903 2148 1937
rect 2114 1835 2148 1869
rect 2900 1808 2934 1842
rect 3087 1808 3121 1842
rect 2900 1740 2934 1774
rect 3087 1740 3121 1774
rect 3258 1808 3292 1842
rect 3258 1740 3292 1774
rect 3559 1808 3593 1842
rect 3559 1740 3593 1774
rect 3730 1808 3764 1842
rect 3730 1740 3764 1774
rect 3912 1808 3946 1842
rect 3912 1740 3946 1774
rect 4083 1808 4117 1842
rect 4083 1740 4117 1774
rect 4387 1808 4421 1842
rect 4387 1740 4421 1774
rect 4558 1808 4592 1842
rect 4558 1740 4592 1774
rect 4861 1808 4895 1842
rect 4861 1740 4895 1774
rect 5039 1808 5073 1842
rect 5039 1740 5073 1774
rect 1558 1227 1592 1261
rect 1634 1227 1668 1261
rect 1711 1227 1745 1261
rect 1788 1227 1822 1261
rect 1904 1227 1938 1261
rect 1972 1227 2006 1261
rect 2262 1227 2296 1261
rect 2338 1227 2372 1261
rect 2415 1227 2449 1261
rect 2492 1227 2526 1261
rect 1525 1022 1559 1056
rect 1601 1022 1635 1056
rect 1678 1022 1712 1056
rect 1755 1022 1789 1056
rect 1871 1022 1905 1056
rect 1939 1022 1973 1056
rect 2229 1022 2263 1056
rect 2305 1022 2339 1056
rect 2382 1022 2416 1056
rect 2459 1022 2493 1056
rect -52 498 -18 532
rect -52 430 -18 464
rect 119 498 153 532
rect 119 430 153 464
rect 421 498 455 532
rect 421 430 455 464
rect 592 498 626 532
rect 779 498 813 532
rect 592 430 626 464
rect 779 430 813 464
rect 1073 498 1107 532
rect 2899 506 2933 540
rect 3086 506 3120 540
rect 1073 430 1107 464
rect 2081 414 2115 448
rect 2081 346 2115 380
rect 2899 438 2933 472
rect 3086 438 3120 472
rect 3258 506 3292 540
rect 3258 438 3292 472
rect 3560 506 3594 540
rect 3560 438 3594 472
rect 3731 506 3765 540
rect 3731 438 3765 472
rect 4035 506 4069 540
rect 4035 438 4069 472
rect 4206 506 4240 540
rect 4206 438 4240 472
rect 4388 506 4422 540
rect 4388 438 4422 472
rect 4559 506 4593 540
rect 4559 438 4593 472
rect 4864 506 4898 540
rect 4864 438 4898 472
rect 5035 506 5069 540
rect 5035 438 5069 472
rect 1519 28 1553 62
rect 1587 28 1621 62
rect 2047 28 2081 62
rect 2115 28 2149 62
rect 2229 28 2263 62
rect 2305 28 2339 62
rect 2382 28 2416 62
rect 2459 28 2493 62
<< locali >>
rect 2067 3677 2119 3711
rect 2153 3677 2253 3711
rect 2287 3677 2311 3711
rect 2067 3603 2140 3677
rect 2067 3569 2106 3603
rect 2067 3554 2140 3569
rect 2067 3497 2106 3554
rect 2067 3486 2140 3497
rect 2067 3452 2106 3486
rect 2067 3436 2140 3452
rect 2282 3554 2316 3570
rect 2282 3486 2316 3520
rect 2179 3358 2195 3392
rect 2229 3358 2245 3392
rect 2179 3324 2245 3358
rect 2179 3290 2195 3324
rect 2229 3290 2245 3324
rect 2106 3239 2140 3240
rect 2040 3224 2140 3239
rect 2040 3190 2106 3224
rect 2040 3156 2140 3190
rect 2040 3116 2106 3156
rect 2040 3088 2140 3116
rect 2040 3044 2106 3088
rect 2040 3006 2140 3044
rect 2040 2972 2106 3006
rect 2040 2962 2140 2972
rect 2040 2928 2106 2962
rect 2040 2894 2140 2928
rect 2040 2860 2106 2894
rect 2040 2826 2140 2860
rect 2040 2792 2106 2826
rect 2040 2655 2140 2792
rect 2282 3224 2316 3452
rect 2282 3156 2316 3190
rect 2282 3088 2316 3122
rect 2282 2962 2316 3054
rect 2282 2894 2316 2928
rect 2282 2826 2316 2860
rect 2282 2774 2316 2792
rect 2040 2621 2099 2655
rect 2133 2621 2183 2655
rect 2217 2621 2266 2655
rect 2300 2621 2324 2655
rect 2040 2587 2324 2621
rect 2040 2553 2099 2587
rect 2133 2553 2183 2587
rect 2217 2553 2266 2587
rect 2300 2553 2324 2587
rect 1536 2221 1552 2255
rect 1586 2221 1620 2255
rect 1654 2221 2080 2255
rect 2114 2221 2148 2255
rect 2182 2221 2198 2255
rect 2246 2221 2262 2255
rect 2296 2221 2338 2255
rect 2372 2221 2415 2255
rect 2449 2221 2492 2255
rect 2526 2221 2542 2255
rect 2784 2251 2804 2285
rect 2838 2251 2840 2285
rect 2874 2251 2876 2285
rect 2942 2251 2948 2285
rect 3010 2251 3020 2285
rect 3078 2251 3092 2285
rect 3146 2251 3164 2285
rect 3214 2251 3236 2285
rect 3282 2251 3308 2285
rect 3350 2251 3380 2285
rect 3418 2251 3452 2285
rect 3486 2251 3520 2285
rect 3558 2251 3588 2285
rect 3630 2251 3656 2285
rect 3702 2251 3714 2285
rect 1497 2167 1531 2183
rect 306 2112 331 2146
rect 365 2112 371 2146
rect 437 2112 439 2146
rect 473 2112 475 2146
rect 541 2112 547 2146
rect 609 2112 619 2146
rect 677 2112 691 2146
rect 745 2112 763 2146
rect 813 2112 835 2146
rect 881 2112 907 2146
rect 949 2112 979 2146
rect 1017 2112 1051 2146
rect 1085 2112 1119 2146
rect 1157 2112 1187 2146
rect 1229 2112 1255 2146
rect 1301 2112 1313 2146
rect 1497 2099 1531 2133
rect -142 2012 -108 2027
rect -142 1944 -108 1955
rect -142 1894 -108 1910
rect 34 2012 68 2028
rect 34 1944 68 1978
rect -70 1816 -54 1850
rect -20 1816 -4 1850
rect -70 1782 -4 1816
rect -70 1748 -54 1782
rect -20 1748 -4 1782
rect 34 1698 68 1910
rect 210 2012 244 2027
rect 210 1944 244 1955
rect 210 1894 244 1910
rect 334 2012 368 2028
rect 334 1944 368 1978
rect 108 1816 124 1850
rect 166 1816 174 1850
rect 108 1782 174 1816
rect 108 1748 124 1782
rect 158 1778 174 1782
rect 166 1748 174 1778
rect 334 1699 368 1910
rect 510 2012 544 2027
rect 510 1944 544 1955
rect 510 1894 544 1910
rect 686 2012 720 2028
rect 686 1944 720 1978
rect -142 1682 -108 1698
rect 34 1682 244 1698
rect 34 1664 210 1682
rect -142 1614 -108 1648
rect -142 1546 -108 1580
rect -142 1420 -108 1512
rect -142 1352 -108 1386
rect -142 1310 -108 1318
rect -142 1238 -108 1250
rect 34 1614 68 1630
rect 34 1546 68 1580
rect 34 1420 68 1512
rect 34 1352 68 1386
rect 34 1284 68 1318
rect 34 1234 68 1250
rect 210 1614 244 1648
rect 367 1682 368 1699
rect 333 1648 334 1665
rect 333 1627 368 1648
rect 367 1614 368 1627
rect 210 1546 244 1580
rect 210 1477 244 1512
rect 210 1420 244 1443
rect 210 1352 244 1371
rect 210 1284 244 1318
rect 210 1204 244 1250
rect 334 1546 368 1580
rect 334 1420 368 1512
rect 334 1352 368 1386
rect 405 1816 421 1850
rect 455 1816 471 1850
rect 405 1782 471 1816
rect 405 1748 421 1782
rect 455 1748 471 1782
rect 576 1816 592 1850
rect 626 1816 642 1850
rect 686 1845 720 1910
rect 862 2012 896 2027
rect 862 1944 896 1955
rect 862 1894 896 1910
rect 1038 2012 1072 2028
rect 1038 1944 1072 1978
rect 576 1782 642 1816
rect 576 1748 592 1782
rect 626 1748 642 1782
rect 405 1484 471 1748
rect 580 1699 642 1748
rect 719 1811 720 1845
rect 685 1773 720 1811
rect 719 1739 720 1773
rect 405 1450 421 1484
rect 455 1450 471 1484
rect 405 1412 471 1450
rect 405 1378 421 1412
rect 455 1378 471 1412
rect 510 1682 544 1698
rect 510 1614 544 1648
rect 510 1546 544 1580
rect 580 1665 589 1699
rect 623 1665 642 1699
rect 580 1627 642 1665
rect 580 1593 589 1627
rect 623 1593 642 1627
rect 580 1575 642 1593
rect 686 1682 720 1739
rect 686 1614 720 1648
rect 510 1420 544 1512
rect 334 1284 368 1318
rect 334 1232 368 1250
rect 510 1352 544 1386
rect 510 1310 544 1318
rect 510 1238 544 1250
rect 686 1546 720 1580
rect 763 1816 779 1850
rect 813 1816 829 1850
rect 763 1782 829 1816
rect 763 1748 779 1782
rect 813 1748 829 1782
rect 934 1820 949 1850
rect 934 1816 950 1820
rect 984 1816 1000 1850
rect 934 1782 1000 1816
rect 934 1748 949 1782
rect 984 1748 1000 1782
rect 763 1696 827 1748
rect 1038 1698 1072 1910
rect 1214 2012 1248 2027
rect 1214 1944 1248 1955
rect 1214 1894 1248 1910
rect 1497 1939 1531 2065
rect 1673 2167 1707 2183
rect 1673 2099 1707 2125
rect 1673 2049 1707 2053
rect 1531 1905 1569 1939
rect 1112 1816 1128 1850
rect 1162 1816 1178 1850
rect 1112 1782 1178 1816
rect 1112 1748 1128 1782
rect 1162 1748 1178 1782
rect 1497 1765 1531 1905
rect 1741 1830 1815 2221
rect 1849 2167 1883 2183
rect 1849 2099 1883 2133
rect 1849 2049 1883 2065
rect 2025 2167 2059 2183
rect 2025 2099 2059 2133
rect 1917 1862 1991 1864
rect 1741 1796 1758 1830
rect 1792 1796 1815 1830
rect 1919 1828 1957 1862
rect 763 1662 783 1696
rect 817 1662 827 1696
rect 763 1624 827 1662
rect 763 1590 783 1624
rect 817 1590 827 1624
rect 763 1575 827 1590
rect 862 1682 896 1698
rect 1038 1682 1248 1698
rect 1038 1664 1214 1682
rect 862 1614 896 1648
rect 686 1420 720 1512
rect 686 1352 720 1386
rect 686 1284 720 1318
rect 686 1232 720 1250
rect 862 1546 896 1580
rect 862 1420 896 1512
rect 862 1352 896 1386
rect 862 1310 896 1318
rect 862 1238 896 1250
rect 1038 1614 1072 1630
rect 1038 1546 1072 1580
rect 1038 1420 1072 1512
rect 1214 1614 1248 1648
rect 1214 1546 1248 1580
rect 1214 1484 1248 1512
rect 1038 1352 1072 1386
rect 1230 1450 1248 1484
rect 1196 1420 1248 1450
rect 1196 1412 1214 1420
rect 1230 1378 1248 1386
rect 1038 1284 1072 1318
rect 1038 1234 1072 1250
rect 1214 1352 1248 1378
rect 1214 1284 1248 1318
rect 1497 1697 1531 1731
rect 1497 1629 1531 1663
rect 1497 1497 1531 1595
rect 1497 1429 1531 1463
rect 1497 1361 1531 1395
rect 1497 1311 1531 1327
rect 1673 1765 1707 1781
rect 1673 1697 1707 1731
rect 1673 1629 1707 1663
rect 1673 1497 1707 1595
rect 1673 1429 1707 1463
rect 1673 1361 1707 1393
rect 1673 1311 1707 1321
rect 1741 1758 1815 1796
rect 1741 1724 1758 1758
rect 1792 1724 1815 1758
rect 1741 1261 1815 1724
rect 1849 1765 1883 1781
rect 1849 1697 1883 1731
rect 1849 1629 1883 1663
rect 1849 1497 1883 1595
rect 1849 1429 1883 1463
rect 1849 1361 1883 1395
rect 1849 1311 1883 1327
rect 1917 1261 1991 1828
rect 2025 1765 2059 2065
rect 2201 2167 2235 2183
rect 2201 2099 2235 2133
rect 2201 2049 2235 2065
rect 2114 1939 2148 1953
rect 2127 1937 2165 1939
rect 2148 1905 2165 1937
rect 2114 1869 2148 1903
rect 2114 1819 2148 1835
rect 2025 1697 2059 1731
rect 2025 1658 2059 1663
rect 2201 1765 2235 1781
rect 2201 1697 2235 1731
rect 2025 1629 2027 1658
rect 2061 1624 2099 1658
rect 2201 1629 2235 1663
rect 2025 1497 2059 1595
rect 2025 1429 2059 1463
rect 2025 1361 2059 1395
rect 2025 1311 2059 1327
rect 2201 1497 2235 1595
rect 2201 1429 2235 1463
rect 2201 1361 2235 1395
rect 2201 1311 2235 1327
rect 2269 1743 2343 2221
rect 2784 2211 3714 2251
rect 2377 2167 2411 2183
rect 2377 2099 2411 2125
rect 2377 2049 2411 2053
rect 2553 2167 2587 2183
rect 2553 2099 2587 2133
rect 2784 2177 2804 2211
rect 2838 2177 2840 2211
rect 2874 2177 2876 2211
rect 2942 2177 2948 2211
rect 3010 2177 3020 2211
rect 3078 2177 3092 2211
rect 3146 2177 3164 2211
rect 3214 2177 3236 2211
rect 3282 2177 3308 2211
rect 3350 2177 3380 2211
rect 3418 2177 3452 2211
rect 3486 2177 3520 2211
rect 3558 2177 3588 2211
rect 3630 2177 3656 2211
rect 3702 2177 3714 2211
rect 2784 2138 3714 2177
rect 2784 2104 2820 2138
rect 2854 2104 2868 2138
rect 2926 2104 2936 2138
rect 2998 2104 3004 2138
rect 3070 2104 3072 2138
rect 3106 2104 3108 2138
rect 3174 2104 3180 2138
rect 3242 2104 3252 2138
rect 3310 2104 3324 2138
rect 3378 2104 3396 2138
rect 3446 2104 3468 2138
rect 3514 2104 3540 2138
rect 3582 2104 3612 2138
rect 3650 2104 3684 2138
rect 3718 2104 3752 2138
rect 3790 2104 3820 2138
rect 3862 2104 3888 2138
rect 3934 2104 3956 2138
rect 4006 2104 4024 2138
rect 4078 2104 4092 2138
rect 4150 2104 4160 2138
rect 4222 2104 4228 2138
rect 4294 2104 4296 2138
rect 4330 2104 4332 2138
rect 4398 2104 4404 2138
rect 4466 2104 4476 2138
rect 4534 2104 4548 2138
rect 4602 2104 4620 2138
rect 4670 2104 4692 2138
rect 4738 2104 4764 2138
rect 4806 2104 4836 2138
rect 4874 2104 4908 2138
rect 4942 2104 4976 2138
rect 5014 2104 5044 2138
rect 5086 2104 5112 2138
rect 5158 2104 5170 2138
rect 2553 1862 2587 2065
rect 2817 2004 2851 2019
rect 2817 1936 2851 1947
rect 2817 1886 2851 1902
rect 2993 2004 3027 2020
rect 2993 1936 3027 1970
rect 2515 1828 2553 1862
rect 2269 1709 2295 1743
rect 2329 1709 2343 1743
rect 2269 1671 2343 1709
rect 2269 1637 2295 1671
rect 2329 1637 2343 1671
rect 2269 1261 2343 1637
rect 2377 1765 2411 1781
rect 2377 1697 2411 1731
rect 2377 1629 2411 1663
rect 2377 1497 2411 1595
rect 2377 1429 2411 1463
rect 2377 1361 2411 1393
rect 2377 1311 2411 1321
rect 2553 1765 2587 1828
rect 2884 1808 2900 1842
rect 2934 1808 2950 1842
rect 2884 1774 2950 1808
rect 2884 1740 2900 1774
rect 2934 1740 2950 1774
rect 2553 1697 2587 1731
rect 2553 1629 2587 1663
rect 2553 1497 2587 1595
rect 2553 1429 2587 1463
rect 2553 1361 2587 1395
rect 2553 1311 2587 1327
rect 2817 1674 2851 1690
rect 2817 1606 2851 1640
rect 2817 1538 2851 1572
rect 2886 1689 2949 1740
rect 2886 1655 2893 1689
rect 2927 1655 2949 1689
rect 2886 1617 2949 1655
rect 2886 1583 2893 1617
rect 2927 1583 2949 1617
rect 2886 1565 2949 1583
rect 2993 1674 3027 1902
rect 3169 2004 3203 2019
rect 3169 1936 3203 1947
rect 3169 1886 3203 1902
rect 3345 2004 3379 2020
rect 3345 1936 3379 1970
rect 3071 1808 3087 1842
rect 3121 1808 3137 1842
rect 3071 1774 3137 1808
rect 3071 1740 3087 1774
rect 3121 1740 3137 1774
rect 3242 1808 3258 1842
rect 3301 1808 3308 1842
rect 3242 1774 3308 1808
rect 3242 1740 3258 1774
rect 3292 1770 3308 1774
rect 3301 1740 3308 1770
rect 2993 1606 3027 1640
rect 2817 1412 2851 1504
rect 2817 1344 2851 1378
rect 2817 1302 2851 1310
rect 1214 1204 1248 1250
rect 1542 1227 1558 1261
rect 1592 1227 1634 1261
rect 1668 1227 1711 1261
rect 1745 1227 1788 1261
rect 1822 1227 1838 1261
rect 1888 1227 1904 1261
rect 1938 1227 1972 1261
rect 2006 1227 2022 1261
rect 2246 1227 2262 1261
rect 2296 1227 2338 1261
rect 2372 1227 2415 1261
rect 2449 1227 2492 1261
rect 2526 1227 2542 1261
rect 2817 1230 2851 1242
rect 2993 1538 3027 1572
rect 3070 1689 3135 1740
rect 3070 1655 3087 1689
rect 3121 1655 3135 1689
rect 3070 1617 3135 1655
rect 3070 1583 3087 1617
rect 3121 1583 3135 1617
rect 3070 1565 3135 1583
rect 3169 1674 3203 1690
rect 3169 1606 3203 1640
rect 2993 1484 3027 1504
rect 2993 1412 3027 1450
rect 2993 1344 3027 1378
rect 2993 1276 3027 1310
rect 2993 1224 3027 1242
rect 3169 1538 3203 1572
rect 3169 1412 3203 1504
rect 3169 1344 3203 1378
rect 3169 1302 3203 1310
rect 3169 1230 3203 1242
rect 3345 1689 3379 1902
rect 3469 2004 3508 2020
rect 3503 1970 3508 2004
rect 3469 1947 3508 1970
rect 3821 2004 3855 2019
rect 4168 2004 4207 2020
rect 4168 1970 4173 2004
rect 4168 1947 4207 1970
rect 3469 1936 3679 1947
rect 3503 1913 3679 1936
rect 3469 1886 3503 1902
rect 3558 1842 3592 1843
rect 3543 1808 3559 1842
rect 3593 1808 3609 1842
rect 3543 1805 3609 1808
rect 3543 1771 3558 1805
rect 3592 1774 3609 1805
rect 3543 1740 3559 1771
rect 3593 1740 3609 1774
rect 3645 1721 3679 1913
rect 3821 1936 3855 1947
rect 3821 1886 3855 1902
rect 3997 1936 4207 1947
rect 3997 1913 4173 1936
rect 3345 1617 3379 1640
rect 3345 1538 3379 1572
rect 3345 1412 3379 1504
rect 3345 1344 3379 1378
rect 3345 1276 3379 1310
rect 3345 1224 3379 1242
rect 3469 1674 3503 1690
rect 3469 1606 3503 1640
rect 3469 1538 3503 1572
rect 3469 1412 3503 1504
rect 3469 1344 3503 1378
rect 3469 1302 3503 1310
rect 3469 1230 3503 1242
rect 3645 1674 3679 1687
rect 3645 1606 3679 1615
rect 3645 1538 3679 1572
rect 3645 1412 3679 1504
rect 3714 1808 3730 1842
rect 3764 1808 3780 1842
rect 3714 1774 3780 1808
rect 3714 1740 3730 1774
rect 3764 1740 3780 1774
rect 3714 1534 3780 1740
rect 3896 1808 3912 1842
rect 3946 1808 3962 1842
rect 3896 1774 3962 1808
rect 3896 1740 3912 1774
rect 3946 1740 3962 1774
rect 3896 1721 3962 1740
rect 3714 1500 3730 1534
rect 3764 1500 3780 1534
rect 3714 1462 3780 1500
rect 3714 1428 3730 1462
rect 3764 1428 3780 1462
rect 3714 1410 3780 1428
rect 3821 1674 3855 1690
rect 3821 1606 3855 1640
rect 3896 1687 3911 1721
rect 3945 1687 3962 1721
rect 3896 1649 3962 1687
rect 3896 1615 3911 1649
rect 3945 1615 3962 1649
rect 3997 1674 4031 1913
rect 4173 1886 4207 1902
rect 4297 2004 4336 2020
rect 4331 1970 4336 2004
rect 4297 1947 4336 1970
rect 4649 2004 4683 2019
rect 4297 1936 4507 1947
rect 4331 1913 4507 1936
rect 4067 1808 4083 1842
rect 4117 1808 4133 1842
rect 4067 1802 4133 1808
rect 4297 1802 4331 1902
rect 4389 1842 4423 1845
rect 4101 1774 4139 1802
rect 4117 1768 4139 1774
rect 4173 1768 4225 1802
rect 4259 1768 4297 1802
rect 4371 1808 4387 1842
rect 4421 1808 4437 1842
rect 4371 1807 4437 1808
rect 4371 1774 4389 1807
rect 4067 1740 4083 1768
rect 4117 1740 4133 1768
rect 4371 1740 4387 1774
rect 4423 1773 4437 1807
rect 4421 1740 4437 1773
rect 3821 1538 3855 1572
rect 3821 1412 3855 1504
rect 3645 1344 3679 1378
rect 3645 1276 3679 1310
rect 3645 1224 3679 1242
rect 3821 1344 3855 1378
rect 3821 1302 3855 1310
rect 3821 1230 3855 1242
rect 3997 1606 4031 1609
rect 3997 1571 4031 1572
rect 3997 1412 4031 1504
rect 3997 1344 4031 1378
rect 3997 1276 4031 1310
rect 3997 1224 4031 1242
rect 4173 1674 4207 1690
rect 4173 1606 4207 1640
rect 4173 1538 4207 1572
rect 4173 1412 4207 1504
rect 4173 1344 4207 1378
rect 4173 1302 4207 1310
rect 4173 1230 4207 1242
rect 4297 1674 4331 1690
rect 4297 1606 4331 1640
rect 4297 1538 4331 1572
rect 4297 1412 4331 1504
rect 4297 1344 4331 1378
rect 4297 1302 4331 1310
rect 4297 1230 4331 1242
rect 4473 1674 4507 1913
rect 4649 1936 4683 1947
rect 4649 1886 4683 1902
rect 4773 2004 4807 2019
rect 4773 1936 4807 1947
rect 4773 1886 4807 1902
rect 4949 2004 4983 2020
rect 4949 1936 4983 1970
rect 4473 1606 4507 1640
rect 4473 1538 4507 1572
rect 4542 1808 4558 1842
rect 4592 1808 4608 1842
rect 4542 1774 4608 1808
rect 4542 1740 4558 1774
rect 4592 1740 4608 1774
rect 4542 1618 4608 1740
rect 4845 1808 4861 1842
rect 4895 1808 4911 1842
rect 4845 1774 4911 1808
rect 4845 1740 4861 1774
rect 4895 1740 4911 1774
rect 4542 1584 4565 1618
rect 4599 1584 4608 1618
rect 4542 1546 4608 1584
rect 4542 1520 4565 1546
rect 4599 1520 4608 1546
rect 4649 1674 4683 1690
rect 4649 1606 4683 1640
rect 4649 1538 4683 1572
rect 4473 1412 4507 1504
rect 4473 1344 4507 1378
rect 4473 1276 4507 1310
rect 4473 1224 4507 1242
rect 4649 1412 4683 1504
rect 4649 1344 4683 1378
rect 4649 1302 4683 1310
rect 4649 1230 4683 1242
rect 4773 1674 4807 1690
rect 4773 1606 4807 1640
rect 4773 1538 4807 1572
rect 4773 1412 4807 1504
rect 4845 1527 4911 1740
rect 4949 1762 4983 1902
rect 5125 2004 5159 2019
rect 5125 1936 5159 1947
rect 5125 1886 5159 1902
rect 5023 1847 5089 1860
rect 5023 1842 5042 1847
rect 5023 1808 5039 1842
rect 5076 1813 5089 1847
rect 5073 1808 5089 1813
rect 5023 1775 5089 1808
rect 5023 1774 5042 1775
rect 5023 1740 5039 1774
rect 5076 1741 5089 1775
rect 5073 1740 5089 1741
rect 4949 1690 4983 1728
rect 4983 1674 5159 1690
rect 4983 1656 5125 1674
rect 4845 1493 4864 1527
rect 4898 1493 4911 1527
rect 4845 1455 4911 1493
rect 4845 1421 4864 1455
rect 4898 1421 4911 1455
rect 4845 1417 4911 1421
rect 4949 1606 4983 1622
rect 4949 1538 4983 1572
rect 4773 1344 4807 1378
rect 4773 1302 4807 1310
rect 4773 1230 4807 1242
rect 4949 1412 4983 1504
rect 4949 1344 4983 1378
rect 4949 1276 4983 1310
rect 4949 1226 4983 1242
rect 5125 1606 5159 1640
rect 5125 1538 5159 1572
rect 5125 1412 5159 1504
rect 5125 1344 5159 1378
rect 5125 1276 5159 1310
rect 5125 1196 5159 1242
rect 353 1123 425 1157
rect 475 1123 493 1157
rect 547 1123 561 1157
rect 619 1123 629 1157
rect 691 1123 697 1157
rect 763 1123 765 1157
rect 799 1123 801 1157
rect 867 1123 873 1157
rect 935 1123 945 1157
rect 1003 1123 1017 1157
rect 1071 1123 1089 1157
rect 1139 1123 1161 1157
rect 1207 1123 1233 1157
rect 1275 1123 1305 1157
rect 1343 1123 1377 1157
rect 1411 1123 1503 1157
rect 1549 1123 1575 1157
rect 1617 1123 1647 1157
rect 1685 1123 1719 1157
rect 1753 1123 1787 1157
rect 1825 1123 1855 1157
rect 1897 1123 1923 1157
rect 1969 1123 1991 1157
rect 2041 1123 2059 1157
rect 2113 1123 2127 1157
rect 2185 1123 2195 1157
rect 2257 1123 2263 1157
rect 2329 1123 2331 1157
rect 2365 1123 2367 1157
rect 2433 1123 2439 1157
rect 2501 1123 2532 1157
rect 2809 1123 2865 1157
rect 2923 1123 2933 1157
rect 2995 1123 3001 1157
rect 3067 1123 3069 1157
rect 3103 1123 3105 1157
rect 3171 1123 3177 1157
rect 3239 1123 3249 1157
rect 3307 1123 3321 1157
rect 3375 1123 3393 1157
rect 3443 1123 3465 1157
rect 3511 1123 3537 1157
rect 3579 1123 3609 1157
rect 3647 1123 3681 1157
rect 3715 1123 3749 1157
rect 3787 1123 3817 1157
rect 3859 1123 3885 1157
rect 3931 1123 3953 1157
rect 4003 1123 4021 1157
rect 4075 1123 4089 1157
rect 4147 1123 4157 1157
rect 4219 1123 4225 1157
rect 4291 1123 4293 1157
rect 4327 1123 4329 1157
rect 4395 1123 4401 1157
rect 4463 1123 4473 1157
rect 4531 1123 4545 1157
rect 4599 1123 4617 1157
rect 4667 1123 4689 1157
rect 4735 1123 4761 1157
rect 4803 1123 4833 1157
rect 4871 1123 4905 1157
rect 4939 1123 4973 1157
rect 5011 1123 5041 1157
rect 5083 1123 5109 1157
rect 5155 1123 5167 1157
rect -142 1030 -108 1042
rect -142 962 -108 970
rect -142 894 -108 928
rect -142 768 -108 860
rect 34 1030 68 1048
rect 34 962 68 996
rect 34 894 68 928
rect 34 768 68 860
rect -142 700 -108 734
rect -142 632 -108 666
rect 64 719 68 734
rect 30 700 68 719
rect 30 681 34 700
rect 64 647 68 666
rect -142 582 -108 598
rect 34 632 68 647
rect -68 499 -56 532
rect -68 498 -52 499
rect -18 498 -2 532
rect -68 464 -2 498
rect -68 461 -52 464
rect -68 430 -56 461
rect -18 430 -2 464
rect -142 370 -108 386
rect 34 359 68 598
rect 210 1030 244 1042
rect 210 962 244 970
rect 210 894 244 928
rect 210 768 244 860
rect 210 700 244 734
rect 334 1030 368 1048
rect 334 962 368 996
rect 334 894 368 928
rect 334 768 368 860
rect 334 700 368 734
rect 210 632 244 666
rect 210 582 244 598
rect 366 655 368 666
rect 332 632 368 655
rect 332 617 334 632
rect 366 583 368 598
rect 103 498 119 532
rect 153 498 169 532
rect 103 464 169 498
rect 103 430 119 464
rect 153 430 169 464
rect -108 336 68 359
rect -142 325 68 336
rect 210 370 244 386
rect 210 325 244 336
rect -142 302 -103 325
rect -108 268 -103 302
rect -142 252 -103 268
rect 210 253 244 268
rect 334 370 368 583
rect 510 1030 544 1042
rect 510 962 544 970
rect 510 894 544 928
rect 686 1030 720 1048
rect 686 962 720 996
rect 686 896 720 928
rect 510 768 544 860
rect 719 894 720 896
rect 685 860 686 862
rect 685 824 720 860
rect 719 790 720 824
rect 510 700 544 734
rect 686 768 720 790
rect 510 632 544 666
rect 510 582 544 598
rect 579 689 642 707
rect 579 655 589 689
rect 623 655 642 689
rect 579 617 642 655
rect 579 583 589 617
rect 623 583 642 617
rect 579 532 642 583
rect 405 492 421 532
rect 455 492 471 532
rect 405 464 471 492
rect 405 430 421 464
rect 455 430 471 464
rect 576 498 592 532
rect 626 498 642 532
rect 576 464 642 498
rect 576 430 592 464
rect 626 430 642 464
rect 686 700 720 734
rect 862 1030 896 1042
rect 862 962 896 970
rect 862 894 896 928
rect 862 768 896 860
rect 686 632 720 666
rect 334 302 368 336
rect 334 252 368 268
rect 510 370 544 386
rect 510 325 544 336
rect 510 253 544 268
rect 686 370 720 598
rect 763 689 827 707
rect 763 655 783 689
rect 817 655 827 689
rect 763 617 827 655
rect 763 583 783 617
rect 817 583 827 617
rect 763 532 827 583
rect 862 700 896 734
rect 862 632 896 666
rect 862 582 896 598
rect 986 1030 1020 1048
rect 986 962 1020 996
rect 986 894 1020 928
rect 986 768 1020 860
rect 986 700 1020 734
rect 1162 1030 1196 1042
rect 1509 1022 1525 1056
rect 1559 1022 1601 1056
rect 1635 1022 1678 1056
rect 1712 1022 1755 1056
rect 1789 1022 1805 1056
rect 1855 1022 1871 1056
rect 1905 1022 1939 1056
rect 1973 1022 1989 1056
rect 2213 1022 2229 1056
rect 2263 1022 2305 1056
rect 2339 1022 2382 1056
rect 2416 1022 2459 1056
rect 2493 1022 2509 1056
rect 2817 1038 2851 1050
rect 1162 962 1196 970
rect 1162 894 1196 928
rect 1162 768 1196 860
rect 1162 700 1196 734
rect 986 632 1020 666
rect 986 574 1020 598
rect 763 498 779 532
rect 813 498 829 532
rect 763 464 829 498
rect 763 430 779 464
rect 813 430 829 464
rect 986 502 1020 540
rect 686 302 720 336
rect 686 252 720 268
rect 862 370 896 386
rect 862 325 896 336
rect 862 253 896 268
rect 986 370 1020 468
rect 1057 651 1075 685
rect 1109 651 1123 685
rect 1057 613 1123 651
rect 1057 579 1075 613
rect 1109 579 1123 613
rect 1162 632 1196 666
rect 1162 582 1196 598
rect 1464 956 1498 972
rect 1464 888 1498 922
rect 1464 820 1498 854
rect 1464 688 1498 786
rect 1464 620 1498 654
rect 1057 532 1123 579
rect 1057 498 1073 532
rect 1107 498 1123 532
rect 1057 464 1123 498
rect 1057 430 1073 464
rect 1107 430 1123 464
rect 1464 552 1498 586
rect 986 302 1020 336
rect 986 252 1020 268
rect 1162 370 1196 386
rect 1162 325 1196 336
rect 1162 253 1196 268
rect 1464 378 1498 518
rect 1640 962 1674 972
rect 1640 890 1674 922
rect 1640 820 1674 854
rect 1640 688 1674 786
rect 1640 620 1674 654
rect 1640 552 1674 586
rect 1640 502 1674 518
rect 1708 722 1782 1022
rect 1708 688 1728 722
rect 1762 688 1782 722
rect 1708 650 1782 688
rect 1708 616 1728 650
rect 1762 616 1782 650
rect 1498 344 1536 378
rect 1464 218 1498 344
rect 317 117 337 151
rect 371 117 373 151
rect 407 117 409 151
rect 475 117 481 151
rect 543 117 553 151
rect 611 117 625 151
rect 679 117 697 151
rect 747 117 769 151
rect 815 117 841 151
rect 883 117 913 151
rect 951 117 985 151
rect 1019 117 1053 151
rect 1091 117 1121 151
rect 1163 117 1189 151
rect 1235 117 1247 151
rect 1464 150 1498 184
rect 1464 100 1498 116
rect 1640 230 1674 234
rect 1640 158 1674 184
rect 1640 100 1674 116
rect 1708 62 1782 616
rect 1816 956 1850 972
rect 1816 888 1850 922
rect 1816 820 1850 854
rect 1816 688 1850 786
rect 1816 620 1850 654
rect 1816 552 1850 586
rect 1816 502 1850 518
rect 1884 455 1958 1022
rect 1886 421 1924 455
rect 1884 419 1958 421
rect 1992 956 2026 972
rect 1992 888 2026 922
rect 1992 820 2026 854
rect 2168 956 2202 972
rect 2168 888 2202 922
rect 2168 820 2202 854
rect 1992 757 1993 786
rect 2027 757 2065 791
rect 1992 688 2026 757
rect 1992 620 2026 654
rect 1992 552 2026 586
rect 1816 218 1850 234
rect 1816 150 1850 184
rect 1816 100 1850 116
rect 1992 218 2026 518
rect 2168 688 2202 786
rect 2168 620 2202 654
rect 2168 552 2202 586
rect 2168 502 2202 518
rect 2081 448 2115 464
rect 2081 380 2115 414
rect 2115 346 2132 378
rect 2094 344 2132 346
rect 2081 330 2115 344
rect 2236 310 2310 1022
rect 2344 962 2378 972
rect 2344 890 2378 922
rect 2344 820 2378 854
rect 2344 688 2378 786
rect 2344 620 2378 654
rect 2344 552 2378 586
rect 2344 502 2378 518
rect 2520 956 2554 972
rect 2520 888 2554 922
rect 2520 820 2554 854
rect 2520 688 2554 786
rect 2520 620 2554 654
rect 2817 970 2851 978
rect 2817 902 2851 936
rect 2817 776 2851 868
rect 2817 708 2851 742
rect 2993 1038 3027 1056
rect 2993 970 3027 1004
rect 2993 902 3027 936
rect 2993 830 3027 868
rect 2993 776 3027 796
rect 2817 640 2851 674
rect 2817 590 2851 606
rect 2887 697 2949 715
rect 2887 663 2893 697
rect 2927 663 2949 697
rect 2887 625 2949 663
rect 2887 591 2893 625
rect 2927 591 2949 625
rect 2520 552 2554 586
rect 2887 540 2949 591
rect 2520 455 2554 518
rect 2482 421 2520 455
rect 2883 506 2899 540
rect 2933 506 2949 540
rect 2883 472 2949 506
rect 2883 438 2899 472
rect 2933 438 2949 472
rect 2993 708 3027 724
rect 3169 1038 3203 1050
rect 3169 970 3203 978
rect 3169 902 3203 936
rect 3169 776 3203 868
rect 3345 1038 3379 1056
rect 3345 970 3379 1004
rect 3345 902 3379 936
rect 2993 640 3027 674
rect 2257 276 2295 310
rect 1992 150 2026 184
rect 1992 100 2026 116
rect 2168 218 2202 234
rect 2168 150 2202 184
rect 2168 100 2202 116
rect 2236 62 2310 276
rect 2344 230 2378 234
rect 2344 158 2378 184
rect 2344 100 2378 116
rect 2520 218 2554 421
rect 2817 378 2851 394
rect 2817 333 2851 344
rect 2817 261 2851 276
rect 2993 378 3027 606
rect 3070 697 3134 715
rect 3070 663 3087 697
rect 3121 663 3134 697
rect 3070 625 3134 663
rect 3070 591 3087 625
rect 3121 591 3134 625
rect 3070 540 3134 591
rect 3169 708 3203 742
rect 3169 640 3203 674
rect 3169 590 3203 606
rect 3242 796 3261 830
rect 3295 796 3308 830
rect 3242 758 3308 796
rect 3242 724 3261 758
rect 3295 724 3308 758
rect 3242 540 3308 724
rect 3070 506 3086 540
rect 3120 506 3136 540
rect 3070 472 3136 506
rect 3070 438 3086 472
rect 3120 438 3136 472
rect 3242 506 3258 540
rect 3292 506 3308 540
rect 3242 472 3308 506
rect 3242 438 3258 472
rect 3292 438 3308 472
rect 3345 776 3379 868
rect 3345 708 3379 742
rect 3345 640 3379 663
rect 2993 310 3027 344
rect 2993 260 3027 276
rect 3169 378 3203 394
rect 3169 333 3203 344
rect 3169 261 3203 276
rect 3345 378 3379 591
rect 3469 1038 3503 1050
rect 3469 970 3503 978
rect 3469 902 3503 936
rect 3469 776 3503 868
rect 3469 708 3503 742
rect 3469 640 3503 674
rect 3469 590 3503 606
rect 3645 1038 3679 1056
rect 3645 970 3679 1004
rect 3645 902 3679 936
rect 3645 837 3679 868
rect 3821 1038 3855 1050
rect 3821 970 3855 978
rect 3821 902 3855 936
rect 3645 776 3679 803
rect 3645 708 3679 731
rect 3645 640 3679 674
rect 3544 521 3559 540
rect 3544 506 3560 521
rect 3594 506 3610 540
rect 3544 483 3610 506
rect 3544 449 3559 483
rect 3593 472 3610 483
rect 3544 438 3560 449
rect 3594 438 3610 472
rect 3345 310 3379 344
rect 3345 260 3379 276
rect 3469 378 3503 394
rect 3469 333 3503 344
rect 3645 367 3679 606
rect 3715 805 3737 837
rect 3771 805 3781 837
rect 3715 767 3781 805
rect 3715 733 3737 767
rect 3771 733 3781 767
rect 3715 540 3781 733
rect 3821 776 3855 868
rect 3821 708 3855 742
rect 3821 640 3855 674
rect 3821 590 3855 606
rect 3945 1038 3979 1050
rect 3945 970 3979 978
rect 3945 902 3979 936
rect 3945 776 3979 868
rect 3945 708 3979 742
rect 3945 640 3979 674
rect 3945 590 3979 606
rect 4121 1038 4155 1056
rect 4121 970 4155 1004
rect 4121 902 4155 936
rect 4121 839 4155 868
rect 4121 776 4155 805
rect 4121 708 4155 733
rect 4121 640 4155 674
rect 3715 506 3731 540
rect 3765 506 3781 540
rect 3715 472 3781 506
rect 3715 438 3731 472
rect 3765 438 3781 472
rect 4019 506 4035 540
rect 4070 521 4085 540
rect 4069 506 4085 521
rect 4019 483 4085 506
rect 4019 472 4036 483
rect 4019 438 4035 472
rect 4070 449 4085 483
rect 4069 438 4085 449
rect 3821 378 3855 394
rect 3645 344 3821 367
rect 3645 333 3855 344
rect 3469 261 3503 276
rect 3816 310 3855 333
rect 3816 276 3821 310
rect 3816 260 3855 276
rect 3945 378 3979 394
rect 4121 367 4155 606
rect 4297 1038 4331 1050
rect 4297 970 4331 978
rect 4297 902 4331 936
rect 4297 776 4331 868
rect 4297 708 4331 742
rect 4297 640 4331 674
rect 4297 590 4331 606
rect 4473 1038 4507 1056
rect 4473 970 4507 1004
rect 4473 902 4507 936
rect 4473 776 4507 868
rect 4473 708 4507 742
rect 4649 1038 4683 1050
rect 4649 970 4683 978
rect 4649 902 4683 936
rect 4649 776 4683 868
rect 4649 708 4683 742
rect 4473 673 4474 674
rect 4473 640 4508 673
rect 4507 635 4508 640
rect 4473 601 4474 606
rect 4649 640 4683 674
rect 4372 540 4392 559
rect 4190 506 4206 540
rect 4243 521 4256 540
rect 4240 506 4256 521
rect 4190 483 4256 506
rect 4190 472 4209 483
rect 4190 438 4206 472
rect 4243 449 4256 483
rect 4240 438 4256 449
rect 4372 506 4388 540
rect 4426 525 4438 559
rect 4422 506 4438 525
rect 4372 487 4438 506
rect 4372 472 4392 487
rect 4372 438 4388 472
rect 4426 453 4438 487
rect 4422 438 4438 453
rect 3979 344 4155 367
rect 3945 333 4155 344
rect 4297 378 4331 394
rect 4297 333 4331 344
rect 4473 367 4507 601
rect 4649 590 4683 606
rect 4773 1038 4807 1050
rect 4773 970 4807 978
rect 4949 1038 4983 1056
rect 4949 970 4983 1004
rect 4773 902 4807 936
rect 4773 776 4807 868
rect 4773 708 4807 742
rect 4773 640 4807 674
rect 4773 590 4807 606
rect 4848 925 4914 937
rect 4848 891 4860 925
rect 4894 891 4914 925
rect 4848 853 4914 891
rect 4848 819 4860 853
rect 4894 819 4914 853
rect 4543 540 4561 559
rect 4543 506 4559 540
rect 4595 525 4609 559
rect 4593 506 4609 525
rect 4543 487 4609 506
rect 4543 472 4561 487
rect 4543 438 4559 472
rect 4595 453 4609 487
rect 4593 438 4609 453
rect 4848 540 4914 819
rect 4848 506 4864 540
rect 4898 506 4914 540
rect 4848 472 4914 506
rect 4848 438 4864 472
rect 4898 438 4914 472
rect 4949 902 4983 936
rect 4949 810 4983 868
rect 4949 738 4983 742
rect 4949 640 4983 674
rect 4649 378 4683 394
rect 4473 344 4649 367
rect 4473 333 4683 344
rect 3945 310 3984 333
rect 3979 276 3984 310
rect 3945 260 3984 276
rect 4297 261 4331 276
rect 4644 310 4683 333
rect 4644 276 4649 310
rect 4644 260 4683 276
rect 4773 378 4807 394
rect 4773 333 4807 344
rect 4949 367 4983 606
rect 5125 1038 5159 1050
rect 5125 970 5159 978
rect 5125 902 5159 936
rect 5125 776 5159 868
rect 5125 708 5159 742
rect 5125 640 5159 674
rect 5125 590 5159 606
rect 5019 528 5033 540
rect 5019 506 5035 528
rect 5069 506 5085 540
rect 5019 490 5085 506
rect 5019 456 5033 490
rect 5067 472 5085 490
rect 5019 438 5035 456
rect 5069 438 5085 472
rect 5125 378 5159 394
rect 4949 344 5125 367
rect 4949 333 5159 344
rect 4773 261 4807 276
rect 5120 310 5159 333
rect 5120 276 5125 310
rect 5120 260 5159 276
rect 2520 150 2554 184
rect 2805 142 2817 176
rect 2851 142 2865 176
rect 2923 142 2933 176
rect 2995 142 3001 176
rect 3067 142 3069 176
rect 3103 142 3105 176
rect 3171 142 3177 176
rect 3239 142 3249 176
rect 3307 142 3321 176
rect 3375 142 3393 176
rect 3443 142 3465 176
rect 3511 142 3537 176
rect 3579 142 3609 176
rect 3647 142 3681 176
rect 3715 142 3749 176
rect 3787 142 3817 176
rect 3859 142 3885 176
rect 3931 142 3953 176
rect 4003 142 4021 176
rect 4075 142 4089 176
rect 4147 142 4157 176
rect 4219 142 4225 176
rect 4291 142 4293 176
rect 4327 142 4329 176
rect 4395 142 4401 176
rect 4463 142 4473 176
rect 4531 142 4545 176
rect 4599 142 4617 176
rect 4667 142 4689 176
rect 4735 142 4761 176
rect 4803 142 4833 176
rect 4871 142 4905 176
rect 4939 142 4973 176
rect 5011 142 5041 176
rect 5083 142 5109 176
rect 5155 142 5167 176
rect 2520 100 2554 116
rect 1503 28 1519 62
rect 1553 28 1587 62
rect 1621 28 2047 62
rect 2081 28 2115 62
rect 2149 28 2165 62
rect 2213 28 2229 62
rect 2263 28 2305 62
rect 2339 28 2382 62
rect 2416 28 2459 62
rect 2493 28 2509 62
<< viali >>
rect 2106 3569 2140 3603
rect 2106 3520 2140 3531
rect 2106 3497 2140 3520
rect 2106 3122 2140 3150
rect 2106 3116 2140 3122
rect 2106 3054 2140 3078
rect 2106 3044 2140 3054
rect 2106 2972 2140 3006
rect 2804 2251 2838 2285
rect 2876 2251 2908 2285
rect 2908 2251 2910 2285
rect 2948 2251 2976 2285
rect 2976 2251 2982 2285
rect 3020 2251 3044 2285
rect 3044 2251 3054 2285
rect 3092 2251 3112 2285
rect 3112 2251 3126 2285
rect 3164 2251 3180 2285
rect 3180 2251 3198 2285
rect 3236 2251 3248 2285
rect 3248 2251 3270 2285
rect 3308 2251 3316 2285
rect 3316 2251 3342 2285
rect 3380 2251 3384 2285
rect 3384 2251 3414 2285
rect 3452 2251 3486 2285
rect 3524 2251 3554 2285
rect 3554 2251 3558 2285
rect 3596 2251 3622 2285
rect 3622 2251 3630 2285
rect 3668 2251 3690 2285
rect 3690 2251 3702 2285
rect 331 2112 365 2146
rect 403 2112 405 2146
rect 405 2112 437 2146
rect 475 2112 507 2146
rect 507 2112 509 2146
rect 547 2112 575 2146
rect 575 2112 581 2146
rect 619 2112 643 2146
rect 643 2112 653 2146
rect 691 2112 711 2146
rect 711 2112 725 2146
rect 763 2112 779 2146
rect 779 2112 797 2146
rect 835 2112 847 2146
rect 847 2112 869 2146
rect 907 2112 915 2146
rect 915 2112 941 2146
rect 979 2112 983 2146
rect 983 2112 1013 2146
rect 1051 2112 1085 2146
rect 1123 2112 1153 2146
rect 1153 2112 1157 2146
rect 1195 2112 1221 2146
rect 1221 2112 1229 2146
rect 1267 2112 1289 2146
rect 1289 2112 1301 2146
rect -142 2027 -108 2061
rect -142 1978 -108 1989
rect -142 1955 -108 1978
rect -54 1816 -20 1850
rect -54 1748 -20 1778
rect -54 1744 -20 1748
rect 210 2027 244 2061
rect 210 1978 244 1989
rect 210 1955 244 1978
rect 132 1816 158 1850
rect 158 1816 166 1850
rect 132 1748 158 1778
rect 158 1748 166 1778
rect 132 1744 166 1748
rect 510 2027 544 2061
rect 510 1978 544 1989
rect 510 1955 544 1978
rect -142 1284 -108 1310
rect -142 1276 -108 1284
rect -142 1204 -108 1238
rect 333 1682 367 1699
rect 333 1665 334 1682
rect 334 1665 367 1682
rect 333 1614 367 1627
rect 333 1593 334 1614
rect 334 1593 367 1614
rect 210 1443 244 1477
rect 210 1386 244 1405
rect 210 1371 244 1386
rect 862 2027 896 2061
rect 862 1978 896 1989
rect 862 1955 896 1978
rect 949 1850 983 1854
rect 685 1811 719 1845
rect 685 1739 719 1773
rect 421 1450 455 1484
rect 421 1378 455 1412
rect 589 1665 623 1699
rect 589 1593 623 1627
rect 510 1284 544 1310
rect 510 1276 544 1284
rect 510 1204 544 1238
rect 949 1820 950 1850
rect 950 1820 983 1850
rect 949 1748 950 1782
rect 950 1748 983 1782
rect 1214 2027 1248 2061
rect 1214 1978 1248 1989
rect 1214 1955 1248 1978
rect 1673 2133 1707 2159
rect 1673 2125 1707 2133
rect 1673 2065 1707 2087
rect 1673 2053 1707 2065
rect 1497 1905 1531 1939
rect 1569 1905 1603 1939
rect 1128 1850 1162 1853
rect 1128 1819 1162 1850
rect 1128 1748 1162 1781
rect 1758 1796 1792 1830
rect 1885 1828 1919 1862
rect 1957 1828 1991 1862
rect 1128 1747 1162 1748
rect 783 1662 817 1696
rect 783 1590 817 1624
rect 862 1284 896 1310
rect 862 1276 896 1284
rect 862 1204 896 1238
rect 1196 1450 1230 1484
rect 1196 1386 1214 1412
rect 1214 1386 1230 1412
rect 1196 1378 1230 1386
rect 1673 1395 1707 1427
rect 1673 1393 1707 1395
rect 1673 1327 1707 1355
rect 1673 1321 1707 1327
rect 1758 1724 1792 1758
rect 2093 1937 2127 1939
rect 2093 1905 2114 1937
rect 2114 1905 2127 1937
rect 2165 1905 2199 1939
rect 2027 1629 2061 1658
rect 2027 1624 2059 1629
rect 2059 1624 2061 1629
rect 2099 1624 2133 1658
rect 2377 2133 2411 2159
rect 2377 2125 2411 2133
rect 2377 2065 2411 2087
rect 2377 2053 2411 2065
rect 2804 2177 2838 2211
rect 2876 2177 2908 2211
rect 2908 2177 2910 2211
rect 2948 2177 2976 2211
rect 2976 2177 2982 2211
rect 3020 2177 3044 2211
rect 3044 2177 3054 2211
rect 3092 2177 3112 2211
rect 3112 2177 3126 2211
rect 3164 2177 3180 2211
rect 3180 2177 3198 2211
rect 3236 2177 3248 2211
rect 3248 2177 3270 2211
rect 3308 2177 3316 2211
rect 3316 2177 3342 2211
rect 3380 2177 3384 2211
rect 3384 2177 3414 2211
rect 3452 2177 3486 2211
rect 3524 2177 3554 2211
rect 3554 2177 3558 2211
rect 3596 2177 3622 2211
rect 3622 2177 3630 2211
rect 3668 2177 3690 2211
rect 3690 2177 3702 2211
rect 2820 2104 2854 2138
rect 2892 2104 2902 2138
rect 2902 2104 2926 2138
rect 2964 2104 2970 2138
rect 2970 2104 2998 2138
rect 3036 2104 3038 2138
rect 3038 2104 3070 2138
rect 3108 2104 3140 2138
rect 3140 2104 3142 2138
rect 3180 2104 3208 2138
rect 3208 2104 3214 2138
rect 3252 2104 3276 2138
rect 3276 2104 3286 2138
rect 3324 2104 3344 2138
rect 3344 2104 3358 2138
rect 3396 2104 3412 2138
rect 3412 2104 3430 2138
rect 3468 2104 3480 2138
rect 3480 2104 3502 2138
rect 3540 2104 3548 2138
rect 3548 2104 3574 2138
rect 3612 2104 3616 2138
rect 3616 2104 3646 2138
rect 3684 2104 3718 2138
rect 3756 2104 3786 2138
rect 3786 2104 3790 2138
rect 3828 2104 3854 2138
rect 3854 2104 3862 2138
rect 3900 2104 3922 2138
rect 3922 2104 3934 2138
rect 3972 2104 3990 2138
rect 3990 2104 4006 2138
rect 4044 2104 4058 2138
rect 4058 2104 4078 2138
rect 4116 2104 4126 2138
rect 4126 2104 4150 2138
rect 4188 2104 4194 2138
rect 4194 2104 4222 2138
rect 4260 2104 4262 2138
rect 4262 2104 4294 2138
rect 4332 2104 4364 2138
rect 4364 2104 4366 2138
rect 4404 2104 4432 2138
rect 4432 2104 4438 2138
rect 4476 2104 4500 2138
rect 4500 2104 4510 2138
rect 4548 2104 4568 2138
rect 4568 2104 4582 2138
rect 4620 2104 4636 2138
rect 4636 2104 4654 2138
rect 4692 2104 4704 2138
rect 4704 2104 4726 2138
rect 4764 2104 4772 2138
rect 4772 2104 4798 2138
rect 4836 2104 4840 2138
rect 4840 2104 4870 2138
rect 4908 2104 4942 2138
rect 4980 2104 5010 2138
rect 5010 2104 5014 2138
rect 5052 2104 5078 2138
rect 5078 2104 5086 2138
rect 5124 2104 5146 2138
rect 5146 2104 5158 2138
rect 2817 2019 2851 2053
rect 2817 1970 2851 1981
rect 2817 1947 2851 1970
rect 2481 1828 2515 1862
rect 2553 1828 2587 1862
rect 2295 1709 2329 1743
rect 2295 1637 2329 1671
rect 2377 1395 2411 1427
rect 2377 1393 2411 1395
rect 2377 1327 2411 1355
rect 2377 1321 2411 1327
rect 2893 1655 2927 1689
rect 2893 1583 2927 1617
rect 3169 2019 3203 2053
rect 3169 1970 3203 1981
rect 3169 1947 3203 1970
rect 3267 1808 3292 1842
rect 3292 1808 3301 1842
rect 3267 1740 3292 1770
rect 3292 1740 3301 1770
rect 2817 1276 2851 1302
rect 2817 1268 2851 1276
rect 2817 1196 2851 1230
rect 3267 1736 3301 1740
rect 3087 1655 3121 1689
rect 3087 1583 3121 1617
rect 2993 1450 3027 1484
rect 2993 1378 3027 1412
rect 3169 1276 3203 1302
rect 3169 1268 3203 1276
rect 3169 1196 3203 1230
rect 3821 2019 3855 2053
rect 3821 1970 3855 1981
rect 3821 1947 3855 1970
rect 3558 1843 3592 1877
rect 3558 1774 3592 1805
rect 3558 1771 3559 1774
rect 3559 1771 3592 1774
rect 3345 1674 3379 1689
rect 3345 1655 3379 1674
rect 3345 1606 3379 1617
rect 3345 1583 3379 1606
rect 3469 1276 3503 1302
rect 3469 1268 3503 1276
rect 3469 1196 3503 1230
rect 3645 1687 3679 1721
rect 3645 1640 3679 1649
rect 3645 1615 3679 1640
rect 3730 1500 3764 1534
rect 3730 1428 3764 1462
rect 3911 1687 3945 1721
rect 3911 1615 3945 1649
rect 4649 2019 4683 2053
rect 4649 1970 4683 1981
rect 4649 1947 4683 1970
rect 4389 1845 4423 1879
rect 4067 1774 4101 1802
rect 4067 1768 4083 1774
rect 4083 1768 4101 1774
rect 4139 1768 4173 1802
rect 4225 1768 4259 1802
rect 4297 1768 4331 1802
rect 4389 1774 4423 1807
rect 4389 1773 4421 1774
rect 4421 1773 4423 1774
rect 3997 1640 4031 1643
rect 3821 1276 3855 1302
rect 3821 1268 3855 1276
rect 3821 1196 3855 1230
rect 3997 1609 4031 1640
rect 3997 1538 4031 1571
rect 3997 1537 4031 1538
rect 4173 1276 4207 1302
rect 4173 1268 4207 1276
rect 4173 1196 4207 1230
rect 4297 1276 4331 1302
rect 4297 1268 4331 1276
rect 4297 1196 4331 1230
rect 4773 2019 4807 2053
rect 4773 1970 4807 1981
rect 4773 1947 4807 1970
rect 4565 1584 4599 1618
rect 4565 1512 4599 1546
rect 4649 1276 4683 1302
rect 4649 1268 4683 1276
rect 4649 1196 4683 1230
rect 5125 2019 5159 2053
rect 5125 1970 5159 1981
rect 5125 1947 5159 1970
rect 4949 1728 4983 1762
rect 5042 1842 5076 1847
rect 5042 1813 5073 1842
rect 5073 1813 5076 1842
rect 5042 1774 5076 1775
rect 5042 1741 5073 1774
rect 5073 1741 5076 1774
rect 4949 1656 4983 1690
rect 4864 1493 4898 1527
rect 4864 1421 4898 1455
rect 4773 1276 4807 1302
rect 4773 1268 4807 1276
rect 4773 1196 4807 1230
rect 441 1123 459 1157
rect 459 1123 475 1157
rect 513 1123 527 1157
rect 527 1123 547 1157
rect 585 1123 595 1157
rect 595 1123 619 1157
rect 657 1123 663 1157
rect 663 1123 691 1157
rect 729 1123 731 1157
rect 731 1123 763 1157
rect 801 1123 833 1157
rect 833 1123 835 1157
rect 873 1123 901 1157
rect 901 1123 907 1157
rect 945 1123 969 1157
rect 969 1123 979 1157
rect 1017 1123 1037 1157
rect 1037 1123 1051 1157
rect 1089 1123 1105 1157
rect 1105 1123 1123 1157
rect 1161 1123 1173 1157
rect 1173 1123 1195 1157
rect 1233 1123 1241 1157
rect 1241 1123 1267 1157
rect 1305 1123 1309 1157
rect 1309 1123 1339 1157
rect 1377 1123 1411 1157
rect 1503 1123 1515 1157
rect 1515 1123 1537 1157
rect 1575 1123 1583 1157
rect 1583 1123 1609 1157
rect 1647 1123 1651 1157
rect 1651 1123 1681 1157
rect 1719 1123 1753 1157
rect 1791 1123 1821 1157
rect 1821 1123 1825 1157
rect 1863 1123 1889 1157
rect 1889 1123 1897 1157
rect 1935 1123 1957 1157
rect 1957 1123 1969 1157
rect 2007 1123 2025 1157
rect 2025 1123 2041 1157
rect 2079 1123 2093 1157
rect 2093 1123 2113 1157
rect 2151 1123 2161 1157
rect 2161 1123 2185 1157
rect 2223 1123 2229 1157
rect 2229 1123 2257 1157
rect 2295 1123 2297 1157
rect 2297 1123 2329 1157
rect 2367 1123 2399 1157
rect 2399 1123 2401 1157
rect 2439 1123 2467 1157
rect 2467 1123 2473 1157
rect 2889 1123 2899 1157
rect 2899 1123 2923 1157
rect 2961 1123 2967 1157
rect 2967 1123 2995 1157
rect 3033 1123 3035 1157
rect 3035 1123 3067 1157
rect 3105 1123 3137 1157
rect 3137 1123 3139 1157
rect 3177 1123 3205 1157
rect 3205 1123 3211 1157
rect 3249 1123 3273 1157
rect 3273 1123 3283 1157
rect 3321 1123 3341 1157
rect 3341 1123 3355 1157
rect 3393 1123 3409 1157
rect 3409 1123 3427 1157
rect 3465 1123 3477 1157
rect 3477 1123 3499 1157
rect 3537 1123 3545 1157
rect 3545 1123 3571 1157
rect 3609 1123 3613 1157
rect 3613 1123 3643 1157
rect 3681 1123 3715 1157
rect 3753 1123 3783 1157
rect 3783 1123 3787 1157
rect 3825 1123 3851 1157
rect 3851 1123 3859 1157
rect 3897 1123 3919 1157
rect 3919 1123 3931 1157
rect 3969 1123 3987 1157
rect 3987 1123 4003 1157
rect 4041 1123 4055 1157
rect 4055 1123 4075 1157
rect 4113 1123 4123 1157
rect 4123 1123 4147 1157
rect 4185 1123 4191 1157
rect 4191 1123 4219 1157
rect 4257 1123 4259 1157
rect 4259 1123 4291 1157
rect 4329 1123 4361 1157
rect 4361 1123 4363 1157
rect 4401 1123 4429 1157
rect 4429 1123 4435 1157
rect 4473 1123 4497 1157
rect 4497 1123 4507 1157
rect 4545 1123 4565 1157
rect 4565 1123 4579 1157
rect 4617 1123 4633 1157
rect 4633 1123 4651 1157
rect 4689 1123 4701 1157
rect 4701 1123 4723 1157
rect 4761 1123 4769 1157
rect 4769 1123 4795 1157
rect 4833 1123 4837 1157
rect 4837 1123 4867 1157
rect 4905 1123 4939 1157
rect 4977 1123 5007 1157
rect 5007 1123 5011 1157
rect 5049 1123 5075 1157
rect 5075 1123 5083 1157
rect 5121 1123 5143 1157
rect 5143 1123 5155 1157
rect -142 1042 -108 1076
rect -142 996 -108 1004
rect -142 970 -108 996
rect 30 734 34 753
rect 34 734 64 753
rect 30 719 64 734
rect 30 666 34 681
rect 34 666 64 681
rect 30 647 64 666
rect -56 532 -22 533
rect -56 499 -52 532
rect -52 499 -22 532
rect -56 430 -52 461
rect -52 430 -22 461
rect -56 427 -22 430
rect 210 1042 244 1076
rect 210 996 244 1004
rect 210 970 244 996
rect 332 666 334 689
rect 334 666 366 689
rect 332 655 366 666
rect 332 598 334 617
rect 334 598 366 617
rect 332 583 366 598
rect 119 532 153 533
rect 119 499 153 532
rect 119 430 153 461
rect 119 427 153 430
rect 210 302 244 325
rect 210 291 244 302
rect 210 219 244 253
rect 510 1042 544 1076
rect 510 996 544 1004
rect 510 970 544 996
rect 685 894 719 896
rect 685 862 686 894
rect 686 862 719 894
rect 685 790 719 824
rect 589 655 623 689
rect 589 583 623 617
rect 421 498 455 526
rect 421 492 455 498
rect 421 430 455 454
rect 862 1042 896 1076
rect 862 996 896 1004
rect 862 970 896 996
rect 421 420 455 430
rect 510 302 544 325
rect 510 291 544 302
rect 510 219 544 253
rect 783 655 817 689
rect 783 583 817 617
rect 1162 1042 1196 1076
rect 2817 1050 2851 1084
rect 1162 996 1196 1004
rect 1162 970 1196 996
rect 986 540 1020 574
rect 986 468 1020 502
rect 862 302 896 325
rect 862 291 896 302
rect 862 219 896 253
rect 1075 651 1109 685
rect 1075 579 1109 613
rect 1162 302 1196 325
rect 1162 291 1196 302
rect 1162 219 1196 253
rect 1640 956 1674 962
rect 1640 928 1674 956
rect 1640 888 1674 890
rect 1640 856 1674 888
rect 1728 688 1762 722
rect 1728 616 1762 650
rect 1464 344 1498 378
rect 1536 344 1570 378
rect 337 117 371 151
rect 409 117 441 151
rect 441 117 443 151
rect 481 117 509 151
rect 509 117 515 151
rect 553 117 577 151
rect 577 117 587 151
rect 625 117 645 151
rect 645 117 659 151
rect 697 117 713 151
rect 713 117 731 151
rect 769 117 781 151
rect 781 117 803 151
rect 841 117 849 151
rect 849 117 875 151
rect 913 117 917 151
rect 917 117 947 151
rect 985 117 1019 151
rect 1057 117 1087 151
rect 1087 117 1091 151
rect 1129 117 1155 151
rect 1155 117 1163 151
rect 1201 117 1223 151
rect 1223 117 1235 151
rect 1640 218 1674 230
rect 1640 196 1674 218
rect 1640 150 1674 158
rect 1640 124 1674 150
rect 1852 421 1886 455
rect 1924 421 1958 455
rect 1993 786 2026 791
rect 2026 786 2027 791
rect 1993 757 2027 786
rect 2065 757 2099 791
rect 2060 346 2081 378
rect 2081 346 2094 378
rect 2060 344 2094 346
rect 2132 344 2166 378
rect 2817 1004 2851 1012
rect 2817 978 2851 1004
rect 2344 956 2378 962
rect 2344 928 2378 956
rect 2344 888 2378 890
rect 2344 856 2378 888
rect 2993 796 3027 830
rect 2993 742 3027 758
rect 2993 724 3027 742
rect 2893 663 2927 697
rect 2893 591 2927 625
rect 2448 421 2482 455
rect 2520 421 2554 455
rect 3169 1050 3203 1084
rect 3169 1004 3203 1012
rect 3169 978 3203 1004
rect 2223 276 2257 310
rect 2295 276 2329 310
rect 2344 218 2378 230
rect 2344 196 2378 218
rect 2344 150 2378 158
rect 2344 124 2378 150
rect 2817 310 2851 333
rect 2817 299 2851 310
rect 2817 227 2851 261
rect 3087 663 3121 697
rect 3087 591 3121 625
rect 3261 796 3295 830
rect 3261 724 3295 758
rect 3345 674 3379 697
rect 3345 663 3379 674
rect 3345 606 3379 625
rect 3345 591 3379 606
rect 3169 310 3203 333
rect 3169 299 3203 310
rect 3169 227 3203 261
rect 3469 1050 3503 1084
rect 3469 1004 3503 1012
rect 3469 978 3503 1004
rect 3821 1050 3855 1084
rect 3821 1004 3855 1012
rect 3821 978 3855 1004
rect 3645 803 3679 837
rect 3645 742 3679 765
rect 3645 731 3679 742
rect 3559 540 3593 555
rect 3559 521 3560 540
rect 3560 521 3593 540
rect 3559 472 3593 483
rect 3559 449 3560 472
rect 3560 449 3593 472
rect 3737 805 3771 839
rect 3737 733 3771 767
rect 3945 1050 3979 1084
rect 3945 1004 3979 1012
rect 3945 978 3979 1004
rect 4121 805 4155 839
rect 4121 742 4155 767
rect 4121 733 4155 742
rect 4036 540 4070 555
rect 4036 521 4069 540
rect 4069 521 4070 540
rect 4036 472 4070 483
rect 4036 449 4069 472
rect 4069 449 4070 472
rect 3469 310 3503 333
rect 3469 299 3503 310
rect 3469 227 3503 261
rect 4297 1050 4331 1084
rect 4297 1004 4331 1012
rect 4297 978 4331 1004
rect 4649 1050 4683 1084
rect 4649 1004 4683 1012
rect 4649 978 4683 1004
rect 4474 674 4507 707
rect 4507 674 4508 707
rect 4474 673 4508 674
rect 4474 606 4507 635
rect 4507 606 4508 635
rect 4474 601 4508 606
rect 4209 540 4243 555
rect 4392 540 4426 559
rect 4209 521 4240 540
rect 4240 521 4243 540
rect 4209 472 4243 483
rect 4209 449 4240 472
rect 4240 449 4243 472
rect 4392 525 4422 540
rect 4422 525 4426 540
rect 4392 472 4426 487
rect 4392 453 4422 472
rect 4422 453 4426 472
rect 4773 1050 4807 1084
rect 4773 1004 4807 1012
rect 4773 978 4807 1004
rect 4860 891 4894 925
rect 4860 819 4894 853
rect 4561 540 4595 559
rect 4561 525 4593 540
rect 4593 525 4595 540
rect 4561 472 4595 487
rect 4561 453 4593 472
rect 4593 453 4595 472
rect 4949 776 4983 810
rect 4949 708 4983 738
rect 4949 704 4983 708
rect 4297 310 4331 333
rect 4297 299 4331 310
rect 4297 227 4331 261
rect 5125 1050 5159 1084
rect 5125 1004 5159 1012
rect 5125 978 5159 1004
rect 5033 540 5067 562
rect 5033 528 5035 540
rect 5035 528 5067 540
rect 5033 472 5067 490
rect 5033 456 5035 472
rect 5035 456 5067 472
rect 4773 310 4807 333
rect 4773 299 4807 310
rect 4773 227 4807 261
rect 2817 142 2851 176
rect 2889 142 2899 176
rect 2899 142 2923 176
rect 2961 142 2967 176
rect 2967 142 2995 176
rect 3033 142 3035 176
rect 3035 142 3067 176
rect 3105 142 3137 176
rect 3137 142 3139 176
rect 3177 142 3205 176
rect 3205 142 3211 176
rect 3249 142 3273 176
rect 3273 142 3283 176
rect 3321 142 3341 176
rect 3341 142 3355 176
rect 3393 142 3409 176
rect 3409 142 3427 176
rect 3465 142 3477 176
rect 3477 142 3499 176
rect 3537 142 3545 176
rect 3545 142 3571 176
rect 3609 142 3613 176
rect 3613 142 3643 176
rect 3681 142 3715 176
rect 3753 142 3783 176
rect 3783 142 3787 176
rect 3825 142 3851 176
rect 3851 142 3859 176
rect 3897 142 3919 176
rect 3919 142 3931 176
rect 3969 142 3987 176
rect 3987 142 4003 176
rect 4041 142 4055 176
rect 4055 142 4075 176
rect 4113 142 4123 176
rect 4123 142 4147 176
rect 4185 142 4191 176
rect 4191 142 4219 176
rect 4257 142 4259 176
rect 4259 142 4291 176
rect 4329 142 4361 176
rect 4361 142 4363 176
rect 4401 142 4429 176
rect 4429 142 4435 176
rect 4473 142 4497 176
rect 4497 142 4507 176
rect 4545 142 4565 176
rect 4565 142 4579 176
rect 4617 142 4633 176
rect 4633 142 4651 176
rect 4689 142 4701 176
rect 4701 142 4723 176
rect 4761 142 4769 176
rect 4769 142 4795 176
rect 4833 142 4837 176
rect 4837 142 4867 176
rect 4905 142 4939 176
rect 4977 142 5007 176
rect 5007 142 5011 176
rect 5049 142 5075 176
rect 5075 142 5083 176
rect 5121 142 5143 176
rect 5143 142 5155 176
<< metal1 >>
rect 2052 3603 2383 3683
rect 2052 3569 2106 3603
rect 2140 3569 2383 3603
rect 2052 3531 2383 3569
rect 2052 3497 2106 3531
rect 2140 3497 2383 3531
rect 2052 3468 2383 3497
rect 2192 3308 2231 3357
tri 2092 3154 2100 3162 se
rect 2100 3154 2147 3162
tri 2147 3154 2155 3162 sw
rect 2051 3150 2325 3154
rect 2051 3116 2106 3150
rect 2140 3116 2325 3150
rect 2051 3078 2325 3116
rect 2051 3044 2106 3078
rect 2140 3044 2325 3078
rect 2051 3006 2325 3044
rect 2051 2972 2106 3006
rect 2140 2972 2325 3006
rect 2051 2960 2325 2972
rect 2700 2797 2706 2849
rect 2758 2797 2777 2849
rect 2829 2797 3932 2849
rect 3984 2797 3996 2849
rect 4048 2797 4054 2849
rect 25 2705 31 2757
rect 83 2705 95 2757
rect 147 2705 2486 2757
rect 2538 2705 2550 2757
rect 2602 2705 2608 2757
rect 123 2613 129 2665
rect 181 2613 193 2665
rect 245 2613 2064 2665
rect 2116 2613 2128 2665
rect 2180 2613 3443 2665
rect 3495 2613 3507 2665
rect 3559 2613 4482 2665
rect 4534 2613 4546 2665
rect 4598 2613 4604 2665
rect -139 2521 -133 2573
rect -81 2521 -69 2573
rect -17 2521 1681 2573
rect 1733 2521 1745 2573
rect 1797 2521 4313 2573
rect 4365 2521 4377 2573
rect 4429 2521 4435 2573
rect 1080 2429 1413 2481
rect 1465 2429 1477 2481
rect 1529 2429 4867 2481
rect 4919 2429 4931 2481
rect 4983 2429 4989 2481
rect 1867 2337 1873 2389
rect 1925 2337 1937 2389
rect 1989 2337 4221 2389
rect 4273 2337 4285 2389
rect 4337 2337 4343 2389
rect 2784 2285 3714 2297
rect 2784 2251 2804 2285
rect 2838 2251 2876 2285
rect 2910 2251 2948 2285
rect 2982 2251 3020 2285
rect 3054 2251 3092 2285
rect 3126 2251 3164 2285
rect 3198 2251 3236 2285
rect 3270 2251 3308 2285
rect 3342 2251 3380 2285
rect 3414 2251 3452 2285
rect 3486 2251 3524 2285
rect 3558 2251 3596 2285
rect 3630 2251 3668 2285
rect 3702 2251 3714 2285
tri 2750 2211 2784 2245 se
rect 2784 2211 3714 2251
tri 2742 2203 2750 2211 se
rect 2750 2203 2804 2211
rect -175 2177 2804 2203
rect 2838 2177 2876 2211
rect 2910 2177 2948 2211
rect 2982 2177 3020 2211
rect 3054 2177 3092 2211
rect 3126 2177 3164 2211
rect 3198 2177 3236 2211
rect 3270 2177 3308 2211
rect 3342 2177 3380 2211
rect 3414 2177 3452 2211
rect 3486 2177 3524 2211
rect 3558 2177 3596 2211
rect 3630 2177 3668 2211
rect 3702 2177 3714 2211
rect -175 2159 3714 2177
rect -175 2146 1673 2159
rect -175 2112 331 2146
rect 365 2112 403 2146
rect 437 2112 475 2146
rect 509 2112 547 2146
rect 581 2112 619 2146
rect 653 2112 691 2146
rect 725 2112 763 2146
rect 797 2112 835 2146
rect 869 2112 907 2146
rect 941 2112 979 2146
rect 1013 2112 1051 2146
rect 1085 2112 1123 2146
rect 1157 2112 1195 2146
rect 1229 2112 1267 2146
rect 1301 2125 1673 2146
rect 1707 2125 2377 2159
rect 2411 2150 3714 2159
tri 3714 2150 3861 2297 sw
rect 2411 2138 5171 2150
rect 2411 2125 2820 2138
rect 1301 2112 2820 2125
rect -175 2104 2820 2112
rect 2854 2104 2892 2138
rect 2926 2104 2964 2138
rect 2998 2104 3036 2138
rect 3070 2104 3108 2138
rect 3142 2104 3180 2138
rect 3214 2104 3252 2138
rect 3286 2104 3324 2138
rect 3358 2104 3396 2138
rect 3430 2104 3468 2138
rect 3502 2104 3540 2138
rect 3574 2104 3612 2138
rect 3646 2104 3684 2138
rect 3718 2104 3756 2138
rect 3790 2104 3828 2138
rect 3862 2104 3900 2138
rect 3934 2104 3972 2138
rect 4006 2104 4044 2138
rect 4078 2104 4116 2138
rect 4150 2104 4188 2138
rect 4222 2104 4260 2138
rect 4294 2104 4332 2138
rect 4366 2104 4404 2138
rect 4438 2104 4476 2138
rect 4510 2104 4548 2138
rect 4582 2104 4620 2138
rect 4654 2104 4692 2138
rect 4726 2104 4764 2138
rect 4798 2104 4836 2138
rect 4870 2104 4908 2138
rect 4942 2104 4980 2138
rect 5014 2104 5052 2138
rect 5086 2104 5124 2138
rect 5158 2104 5171 2138
rect -175 2087 5171 2104
tri 5341 2097 5375 2131 nw
rect -175 2061 1673 2087
rect -175 2027 -142 2061
rect -108 2027 210 2061
rect 244 2027 510 2061
rect 544 2027 862 2061
rect 896 2027 1214 2061
rect 1248 2053 1673 2061
rect 1707 2053 2377 2087
rect 2411 2053 5171 2087
rect 1248 2040 2817 2053
rect 1248 2027 1297 2040
rect -175 2019 1297 2027
tri 1297 2019 1318 2040 nw
tri 2742 2019 2763 2040 ne
rect 2763 2019 2817 2040
rect 2851 2019 3169 2053
rect 3203 2019 3821 2053
rect 3855 2019 4649 2053
rect 4683 2019 4773 2053
rect 4807 2019 5125 2053
rect 5159 2019 5171 2053
rect -175 1989 1260 2019
rect -175 1955 -142 1989
rect -108 1955 210 1989
rect 244 1955 510 1989
rect 544 1955 862 1989
rect 896 1955 1214 1989
rect 1248 1955 1260 1989
tri 1260 1982 1297 2019 nw
tri 2763 1998 2784 2019 ne
rect -175 1943 1260 1955
rect 2784 1981 5171 2019
rect 2784 1947 2817 1981
rect 2851 1947 3169 1981
rect 3203 1947 3821 1981
rect 3855 1947 4649 1981
rect 4683 1947 4773 1981
rect 4807 1947 5125 1981
rect 5159 1947 5171 1981
rect 1485 1939 2211 1945
rect 1485 1905 1497 1939
rect 1531 1905 1569 1939
rect 1603 1905 2093 1939
rect 2127 1905 2165 1939
rect 2199 1905 2211 1939
rect 2784 1935 5171 1947
rect 1485 1899 2211 1905
rect 3630 1898 3682 1904
rect 3466 1881 3598 1893
rect -63 1856 -11 1862
rect -63 1792 -11 1804
rect -63 1732 -11 1740
rect 123 1856 175 1862
rect 123 1792 175 1804
rect 123 1732 175 1740
rect 679 1845 756 1857
rect 679 1811 685 1845
rect 719 1811 756 1845
rect 679 1773 756 1811
rect 679 1739 685 1773
rect 719 1739 756 1773
rect 679 1727 756 1739
rect 943 1854 989 1866
rect 943 1820 949 1854
rect 983 1820 989 1854
rect 943 1782 989 1820
rect 943 1748 949 1782
rect 983 1748 989 1782
rect 943 1727 989 1748
rect 1122 1854 1168 1865
rect 1873 1862 2599 1868
tri 1168 1854 1173 1859 sw
rect 1122 1853 1173 1854
rect 1122 1819 1128 1853
rect 1162 1842 1173 1853
tri 1173 1842 1185 1854 sw
rect 1162 1839 1185 1842
tri 1185 1839 1188 1842 sw
rect 1162 1830 1188 1839
tri 1188 1830 1197 1839 sw
rect 1585 1833 1637 1839
rect 1162 1819 1197 1830
tri 1197 1819 1208 1830 sw
rect 1122 1796 1208 1819
tri 1208 1796 1231 1819 sw
tri 1562 1796 1585 1819 se
rect 1122 1794 1231 1796
tri 1231 1794 1233 1796 sw
tri 1560 1794 1562 1796 se
rect 1562 1794 1585 1796
rect 1122 1781 1585 1794
rect 1122 1747 1128 1781
rect 1162 1769 1637 1781
rect 1162 1756 1585 1769
rect 1162 1747 1168 1756
tri 1168 1753 1171 1756 nw
tri 1541 1753 1544 1756 ne
rect 1544 1753 1585 1756
rect 1122 1735 1168 1747
tri 1544 1735 1562 1753 ne
rect 1562 1735 1585 1753
tri 1562 1729 1568 1735 ne
rect 1568 1729 1585 1735
tri 989 1727 991 1729 sw
tri 1568 1727 1570 1729 ne
rect 1570 1727 1585 1729
rect 943 1724 991 1727
tri 991 1724 994 1727 sw
tri 1570 1724 1573 1727 ne
rect 1573 1724 1585 1727
rect 943 1711 994 1724
tri 994 1711 1007 1724 sw
tri 1573 1712 1585 1724 ne
rect 1585 1711 1637 1717
rect 1752 1830 1798 1842
rect 1752 1796 1758 1830
rect 1792 1796 1798 1830
rect 1873 1828 1885 1862
rect 1919 1828 1957 1862
rect 1991 1828 2481 1862
rect 2515 1828 2553 1862
rect 2587 1828 2599 1862
rect 1873 1822 2599 1828
rect 3257 1848 3309 1854
rect 1752 1771 1798 1796
tri 1798 1771 1825 1798 sw
rect 3257 1777 3309 1796
rect 1752 1770 1825 1771
tri 1825 1770 1826 1771 sw
rect 1752 1764 1826 1770
tri 1826 1764 1832 1770 sw
rect 1752 1758 2048 1764
rect 1752 1724 1758 1758
rect 1792 1724 2048 1758
rect 1752 1712 2048 1724
rect 2100 1712 2112 1764
rect 2164 1712 2170 1764
rect 2289 1753 2335 1755
tri 2335 1753 2337 1755 sw
rect 2289 1743 2337 1753
rect 327 1699 373 1711
tri 581 1709 583 1711 se
rect 583 1709 629 1711
tri 629 1709 631 1711 sw
rect 943 1709 1007 1711
tri 1007 1709 1009 1711 sw
rect 2289 1709 2295 1743
rect 2329 1736 2337 1743
tri 2337 1736 2354 1753 sw
tri 2507 1736 2524 1753 se
rect 2524 1747 2576 1753
rect 2329 1732 2354 1736
tri 2354 1732 2358 1736 sw
tri 2503 1732 2507 1736 se
rect 2507 1732 2524 1736
rect 2329 1709 2524 1732
tri 577 1705 581 1709 se
rect 581 1708 631 1709
tri 631 1708 632 1709 sw
rect 943 1708 1009 1709
tri 1009 1708 1010 1709 sw
rect 581 1706 632 1708
tri 632 1706 634 1708 sw
rect 581 1705 634 1706
tri 373 1699 379 1705 sw
tri 571 1699 577 1705 se
rect 577 1699 634 1705
rect 327 1665 333 1699
rect 367 1672 379 1699
tri 379 1672 406 1699 sw
tri 544 1672 571 1699 se
rect 571 1672 589 1699
rect 367 1665 589 1672
rect 623 1696 634 1699
tri 634 1696 644 1706 sw
tri 767 1696 777 1706 se
rect 777 1696 823 1708
rect 623 1672 644 1696
tri 644 1672 668 1696 sw
tri 743 1672 767 1696 se
rect 767 1672 783 1696
rect 623 1665 783 1672
rect 327 1662 783 1665
rect 817 1662 823 1696
rect 327 1627 823 1662
rect 327 1593 333 1627
rect 367 1608 589 1627
rect 367 1593 385 1608
tri 385 1593 400 1608 nw
tri 556 1593 571 1608 ne
rect 571 1593 589 1608
rect 623 1624 823 1627
rect 943 1689 1010 1708
tri 1010 1689 1029 1708 sw
rect 2289 1695 2524 1709
rect 3518 1877 3598 1881
rect 3518 1843 3558 1877
rect 3592 1843 3598 1877
rect 3518 1829 3598 1843
rect 3466 1817 3598 1829
rect 3518 1805 3598 1817
rect 3518 1771 3558 1805
rect 3592 1771 3598 1805
tri 3682 1891 3695 1904 sw
rect 3682 1882 3695 1891
tri 3695 1882 3704 1891 sw
tri 4374 1882 4383 1891 se
rect 4383 1885 4519 1891
rect 4383 1882 4467 1885
rect 3682 1879 4467 1882
rect 3682 1846 4389 1879
rect 3630 1845 4389 1846
rect 4423 1845 4467 1879
rect 3630 1836 4467 1845
rect 3630 1834 3699 1836
rect 3682 1813 3699 1834
tri 3699 1813 3722 1836 nw
tri 4355 1813 4378 1836 ne
rect 4378 1833 4467 1836
rect 4378 1819 4519 1833
rect 4378 1813 4467 1819
rect 3682 1807 3693 1813
tri 3693 1807 3699 1813 nw
tri 4378 1808 4383 1813 ne
rect 3682 1802 3688 1807
tri 3688 1802 3693 1807 nw
rect 4055 1802 4343 1808
tri 3682 1796 3688 1802 nw
rect 3630 1776 3682 1782
rect 3518 1765 3598 1771
rect 3466 1759 3598 1765
rect 4055 1768 4067 1802
rect 4101 1768 4139 1802
rect 4173 1768 4225 1802
rect 4259 1768 4297 1802
rect 4331 1768 4343 1802
rect 4055 1762 4343 1768
rect 4383 1807 4467 1813
rect 4383 1773 4389 1807
rect 4423 1773 4467 1807
rect 4383 1767 4467 1773
rect 4383 1761 4519 1767
rect 4803 1847 5082 1859
rect 4803 1813 5042 1847
rect 5076 1813 5082 1847
tri 4802 1761 4803 1762 se
rect 4803 1761 4862 1813
tri 4862 1779 4896 1813 nw
tri 5002 1779 5036 1813 ne
rect 5036 1775 5082 1813
rect 5540 1805 5851 2006
tri 4800 1759 4802 1761 se
rect 4802 1759 4862 1761
tri 4775 1734 4800 1759 se
rect 4800 1734 4862 1759
rect 3257 1719 3309 1725
rect 3639 1721 3685 1733
tri 3685 1721 3689 1725 sw
tri 3901 1721 3905 1725 se
rect 3905 1721 3951 1733
rect 943 1671 1029 1689
tri 1029 1671 1047 1689 sw
rect 2289 1683 2576 1695
rect 2289 1680 2524 1683
rect 2289 1671 2365 1680
rect 943 1664 1047 1671
tri 1047 1664 1054 1671 sw
rect 943 1658 2145 1664
rect 943 1654 2027 1658
tri 943 1624 973 1654 ne
rect 973 1624 2027 1654
rect 2061 1624 2099 1658
rect 2133 1624 2145 1658
rect 2289 1637 2295 1671
rect 2329 1655 2365 1671
tri 2365 1655 2390 1680 nw
tri 2490 1655 2515 1680 ne
rect 2515 1655 2524 1680
rect 2329 1649 2359 1655
tri 2359 1649 2365 1655 nw
tri 2515 1649 2521 1655 ne
rect 2521 1649 2524 1655
rect 2329 1637 2335 1649
rect 2289 1625 2335 1637
tri 2335 1625 2359 1649 nw
tri 2521 1646 2524 1649 ne
rect 2524 1625 2576 1631
rect 2887 1689 2933 1701
tri 2933 1689 2940 1696 sw
tri 3074 1689 3081 1696 se
rect 3081 1689 3127 1701
tri 3127 1689 3134 1696 sw
tri 3332 1689 3339 1696 se
rect 3339 1689 3385 1701
rect 2887 1655 2893 1689
rect 2927 1662 2940 1689
tri 2940 1662 2967 1689 sw
tri 3047 1662 3074 1689 se
rect 3074 1662 3087 1689
rect 2927 1655 3087 1662
rect 3121 1662 3134 1689
tri 3134 1662 3161 1689 sw
tri 3305 1662 3332 1689 se
rect 3332 1662 3345 1689
rect 3121 1655 3345 1662
rect 3379 1655 3385 1689
rect 623 1608 783 1624
rect 623 1593 638 1608
rect 327 1590 382 1593
tri 382 1590 385 1593 nw
tri 571 1590 574 1593 ne
rect 574 1590 638 1593
tri 638 1590 656 1608 nw
tri 751 1590 769 1608 ne
rect 769 1590 783 1608
rect 817 1590 823 1624
tri 973 1618 979 1624 ne
rect 979 1618 2145 1624
rect 327 1583 375 1590
tri 375 1583 382 1590 nw
tri 574 1583 581 1590 ne
rect 581 1583 631 1590
tri 631 1583 638 1590 nw
tri 769 1583 776 1590 ne
rect 776 1583 823 1590
rect 327 1581 373 1583
tri 373 1581 375 1583 nw
tri 581 1581 583 1583 ne
rect 583 1581 629 1583
tri 629 1581 631 1583 nw
tri 776 1582 777 1583 ne
rect 777 1578 823 1583
rect 2887 1617 3385 1655
rect 2887 1583 2893 1617
rect 2927 1598 3087 1617
rect 2927 1583 2945 1598
tri 2945 1583 2960 1598 nw
tri 3054 1583 3069 1598 ne
rect 3069 1583 3087 1598
rect 3121 1598 3345 1617
rect 3121 1583 3139 1598
tri 3139 1583 3154 1598 nw
tri 3312 1583 3327 1598 ne
rect 3327 1583 3345 1598
rect 3379 1583 3385 1617
rect 3639 1687 3645 1721
rect 3679 1691 3689 1721
tri 3689 1691 3719 1721 sw
tri 3871 1691 3901 1721 se
rect 3901 1691 3911 1721
rect 3679 1687 3911 1691
rect 3945 1687 3951 1721
rect 3639 1649 3951 1687
rect 4095 1682 4101 1734
rect 4153 1682 4165 1734
rect 4217 1728 4241 1734
tri 4241 1728 4247 1734 sw
tri 4769 1728 4775 1734 se
rect 4775 1728 4862 1734
rect 4217 1682 4862 1728
rect 4943 1762 4989 1774
rect 4943 1728 4949 1762
rect 4983 1728 4989 1762
rect 5036 1741 5042 1775
rect 5076 1741 5082 1775
rect 5036 1729 5082 1741
rect 4943 1690 4989 1728
tri 4935 1656 4943 1664 se
rect 4943 1656 4949 1690
rect 4983 1656 4989 1690
rect 7159 1677 7237 1745
tri 4934 1655 4935 1656 se
rect 4935 1655 4989 1656
rect 3639 1615 3645 1649
rect 3679 1645 3911 1649
rect 3679 1640 3714 1645
tri 3714 1640 3719 1645 nw
tri 3871 1640 3876 1645 ne
rect 3876 1640 3911 1645
rect 3679 1625 3699 1640
tri 3699 1625 3714 1640 nw
tri 3876 1625 3891 1640 ne
rect 3891 1625 3911 1640
rect 3679 1618 3692 1625
tri 3692 1618 3699 1625 nw
tri 3891 1618 3898 1625 ne
rect 3898 1618 3911 1625
rect 3679 1615 3689 1618
tri 3689 1615 3692 1618 nw
tri 3898 1615 3901 1618 ne
rect 3901 1615 3911 1618
rect 3945 1615 3951 1649
rect 3639 1603 3685 1615
tri 3685 1611 3689 1615 nw
tri 3901 1611 3905 1615 ne
rect 3905 1603 3951 1615
rect 3984 1649 4037 1655
rect 2887 1571 2933 1583
tri 2933 1571 2945 1583 nw
tri 3069 1571 3081 1583 ne
rect 3081 1571 3127 1583
tri 3127 1571 3139 1583 nw
tri 3327 1571 3339 1583 ne
rect 3339 1571 3385 1583
rect 4036 1597 4037 1649
tri 4925 1646 4934 1655 se
rect 4934 1646 4989 1655
tri 4919 1640 4925 1646 se
rect 4925 1640 4989 1646
rect 3984 1583 4037 1597
rect 3724 1534 3770 1546
rect 3724 1500 3730 1534
rect 3764 1500 3770 1534
rect 4036 1531 4037 1583
rect 3984 1525 4037 1531
rect 4200 1634 4252 1640
tri 4252 1630 4262 1640 sw
tri 4909 1630 4919 1640 se
rect 4919 1630 4989 1640
rect 4252 1625 4262 1630
tri 4262 1625 4267 1630 sw
rect 4252 1624 4267 1625
tri 4267 1624 4268 1625 sw
rect 4252 1582 4520 1624
rect 4200 1578 4520 1582
rect 4200 1570 4252 1578
tri 4252 1552 4278 1578 nw
tri 4440 1552 4466 1578 ne
rect 4466 1552 4520 1578
tri 4466 1550 4468 1552 ne
rect 4468 1550 4520 1552
rect 4200 1512 4252 1518
rect 4291 1544 4343 1550
tri 4468 1546 4472 1550 ne
rect 4472 1546 4520 1550
tri 4472 1544 4474 1546 ne
rect 3724 1499 3770 1500
tri 3770 1499 3779 1508 sw
tri 4282 1499 4291 1508 se
rect 410 1493 462 1499
rect 3724 1496 3779 1499
tri 3779 1496 3782 1499 sw
tri 4279 1496 4282 1499 se
rect 4282 1496 4291 1499
rect 201 1483 253 1489
rect 201 1417 253 1431
tri 462 1484 466 1488 sw
tri 1186 1484 1190 1488 se
rect 1190 1484 1236 1496
rect 462 1454 466 1484
tri 466 1454 496 1484 sw
tri 1156 1454 1186 1484 se
rect 1186 1454 1196 1484
rect 462 1450 1196 1454
rect 1230 1450 1236 1484
rect 462 1441 1236 1450
rect 410 1424 1236 1441
rect 2987 1484 3033 1496
rect 2987 1450 2993 1484
rect 3027 1450 3033 1484
tri 1656 1428 1667 1439 se
rect 1667 1428 2417 1439
tri 2417 1428 2428 1439 sw
tri 1655 1427 1656 1428 se
rect 1656 1427 2428 1428
rect 462 1412 1236 1424
rect 462 1408 1196 1412
rect 462 1378 466 1408
tri 466 1378 496 1408 nw
tri 1156 1378 1186 1408 ne
rect 1186 1378 1196 1408
rect 1230 1378 1236 1412
tri 1621 1393 1655 1427 se
rect 1655 1393 1673 1427
rect 1707 1393 2377 1427
rect 2411 1421 2428 1427
tri 2428 1421 2435 1428 sw
rect 2411 1418 2435 1421
tri 2435 1418 2438 1421 sw
rect 2411 1412 2438 1418
tri 2438 1412 2444 1418 sw
rect 2987 1412 3033 1450
rect 3724 1493 3782 1496
tri 3782 1493 3785 1496 sw
tri 4276 1493 4279 1496 se
rect 4279 1493 4291 1496
rect 3724 1474 3785 1493
tri 3785 1474 3804 1493 sw
tri 4257 1474 4276 1493 se
rect 4276 1492 4291 1493
rect 4276 1480 4343 1492
rect 4276 1474 4291 1480
rect 3724 1462 4291 1474
rect 3724 1428 3730 1462
rect 3764 1428 4291 1462
rect 3724 1422 4343 1428
rect 4474 1496 4520 1546
rect 4559 1618 4989 1630
tri 7077 1625 7098 1646 ne
rect 7098 1625 7332 1646
tri 7098 1618 7105 1625 ne
rect 7105 1618 7332 1625
rect 4559 1584 4565 1618
rect 4599 1584 4989 1618
tri 7105 1616 7107 1618 ne
rect 7107 1616 7332 1618
tri 7332 1616 7362 1646 nw
rect 4559 1578 4633 1584
tri 4633 1578 4639 1584 nw
rect 4559 1546 4605 1578
tri 4605 1550 4633 1578 nw
rect 4559 1512 4565 1546
rect 4599 1512 4605 1546
rect 7159 1541 7237 1609
rect 4559 1500 4605 1512
rect 4858 1527 4904 1539
tri 4520 1496 4522 1498 sw
tri 4856 1496 4858 1498 se
rect 4858 1496 4864 1527
rect 4474 1493 4522 1496
tri 4522 1493 4525 1496 sw
tri 4853 1493 4856 1496 se
rect 4856 1493 4864 1496
rect 4898 1493 4904 1527
rect 4474 1490 4525 1493
tri 4525 1490 4528 1493 sw
tri 4850 1490 4853 1493 se
rect 4853 1490 4904 1493
tri 5341 1490 5375 1524 sw
rect 4474 1464 4528 1490
tri 4528 1464 4554 1490 sw
tri 4824 1464 4850 1490 se
rect 4850 1464 4904 1490
rect 4474 1455 4904 1464
rect 3724 1421 3775 1422
tri 3775 1421 3776 1422 nw
rect 4474 1421 4864 1455
rect 4898 1421 4904 1455
rect 5798 1449 5833 1488
rect 6826 1452 6865 1496
rect 3724 1418 3772 1421
tri 3772 1418 3775 1421 nw
rect 4474 1418 4904 1421
rect 3724 1416 3770 1418
tri 3770 1416 3772 1418 nw
tri 4673 1416 4675 1418 ne
rect 4675 1416 4808 1418
tri 4675 1412 4679 1416 ne
rect 4679 1412 4808 1416
tri 4808 1412 4814 1418 nw
tri 4849 1412 4855 1418 ne
rect 4855 1412 4904 1418
rect 2411 1409 2444 1412
tri 2444 1409 2447 1412 sw
rect 2411 1393 2447 1409
tri 1606 1378 1621 1393 se
rect 1621 1378 2447 1393
tri 2447 1378 2478 1409 sw
rect 2987 1378 2993 1412
rect 3027 1378 3033 1412
tri 4855 1409 4858 1412 ne
rect 4858 1409 4904 1412
rect 7371 1409 7459 1454
tri 462 1374 466 1378 nw
tri 1186 1374 1190 1378 ne
rect 410 1366 462 1372
rect 1190 1366 1236 1378
tri 1594 1366 1606 1378 se
rect 1606 1366 2478 1378
tri 2478 1366 2490 1378 sw
rect 2987 1366 3033 1378
rect 201 1359 253 1365
tri 1587 1359 1594 1366 se
rect 1594 1359 2490 1366
tri 2490 1359 2497 1366 sw
tri 1583 1355 1587 1359 se
rect 1587 1355 2497 1359
tri 1551 1323 1583 1355 se
rect 1583 1323 1673 1355
rect -154 1321 1673 1323
rect 1707 1321 2377 1355
rect 2411 1323 2497 1355
tri 2497 1323 2533 1359 sw
rect 2411 1321 2533 1323
rect -154 1315 2533 1321
tri 2533 1315 2541 1323 sw
rect -154 1310 5171 1315
rect -154 1276 -142 1310
rect -108 1276 510 1310
rect 544 1276 862 1310
rect 896 1302 5171 1310
rect 896 1276 2817 1302
rect -154 1268 2817 1276
rect 2851 1268 3169 1302
rect 3203 1268 3469 1302
rect 3503 1268 3821 1302
rect 3855 1268 4173 1302
rect 4207 1268 4297 1302
rect 4331 1268 4649 1302
rect 4683 1268 4773 1302
rect 4807 1268 5171 1302
rect -154 1238 5171 1268
rect -154 1204 -142 1238
rect -108 1204 510 1238
rect 544 1204 862 1238
rect 896 1230 5171 1238
rect 896 1204 2817 1230
rect -154 1196 2817 1204
rect 2851 1196 3169 1230
rect 3203 1196 3469 1230
rect 3503 1196 3821 1230
rect 3855 1196 4173 1230
rect 4207 1196 4297 1230
rect 4331 1196 4649 1230
rect 4683 1196 4773 1230
rect 4807 1196 5171 1230
tri -185 1160 -154 1191 se
rect -154 1168 5171 1196
tri 5171 1168 5202 1199 sw
rect -154 1160 5202 1168
rect -185 1157 5202 1160
rect -185 1123 441 1157
rect 475 1123 513 1157
rect 547 1123 585 1157
rect 619 1123 657 1157
rect 691 1123 729 1157
rect 763 1123 801 1157
rect 835 1123 873 1157
rect 907 1123 945 1157
rect 979 1123 1017 1157
rect 1051 1123 1089 1157
rect 1123 1123 1161 1157
rect 1195 1123 1233 1157
rect 1267 1123 1305 1157
rect 1339 1123 1377 1157
rect 1411 1123 1503 1157
rect 1537 1123 1575 1157
rect 1609 1123 1647 1157
rect 1681 1123 1719 1157
rect 1753 1123 1791 1157
rect 1825 1123 1863 1157
rect 1897 1123 1935 1157
rect 1969 1123 2007 1157
rect 2041 1123 2079 1157
rect 2113 1123 2151 1157
rect 2185 1123 2223 1157
rect 2257 1123 2295 1157
rect 2329 1123 2367 1157
rect 2401 1123 2439 1157
rect 2473 1123 2889 1157
rect 2923 1123 2961 1157
rect 2995 1123 3033 1157
rect 3067 1123 3105 1157
rect 3139 1123 3177 1157
rect 3211 1123 3249 1157
rect 3283 1123 3321 1157
rect 3355 1123 3393 1157
rect 3427 1123 3465 1157
rect 3499 1123 3537 1157
rect 3571 1123 3609 1157
rect 3643 1123 3681 1157
rect 3715 1123 3753 1157
rect 3787 1123 3825 1157
rect 3859 1123 3897 1157
rect 3931 1123 3969 1157
rect 4003 1123 4041 1157
rect 4075 1123 4113 1157
rect 4147 1123 4185 1157
rect 4219 1123 4257 1157
rect 4291 1123 4329 1157
rect 4363 1123 4401 1157
rect 4435 1123 4473 1157
rect 4507 1123 4545 1157
rect 4579 1123 4617 1157
rect 4651 1123 4689 1157
rect 4723 1123 4761 1157
rect 4795 1123 4833 1157
rect 4867 1123 4905 1157
rect 4939 1123 4977 1157
rect 5011 1123 5049 1157
rect 5083 1123 5121 1157
rect 5155 1123 5202 1157
rect 5483 1123 5522 1168
rect -185 1084 5202 1123
rect -185 1076 2817 1084
rect -185 1042 -142 1076
rect -108 1042 210 1076
rect 244 1042 510 1076
rect 544 1042 862 1076
rect 896 1042 1162 1076
rect 1196 1050 2817 1076
rect 2851 1050 3169 1084
rect 3203 1050 3469 1084
rect 3503 1050 3821 1084
rect 3855 1050 3945 1084
rect 3979 1050 4297 1084
rect 4331 1050 4649 1084
rect 4683 1050 4773 1084
rect 4807 1050 5125 1084
rect 5159 1050 5202 1084
rect 1196 1042 5202 1050
rect -185 1012 5202 1042
rect -185 1004 2817 1012
rect -185 970 -142 1004
rect -108 970 210 1004
rect 244 970 510 1004
rect 544 970 862 1004
rect 896 970 1162 1004
rect 1196 978 2817 1004
rect 2851 978 3169 1012
rect 3203 978 3469 1012
rect 3503 978 3821 1012
rect 3855 978 3945 1012
rect 3979 978 4297 1012
rect 4331 978 4649 1012
rect 4683 978 4773 1012
rect 4807 978 5125 1012
rect 5159 978 5202 1012
rect 1196 970 5202 978
rect -185 965 5202 970
rect -185 962 2497 965
rect -185 957 1640 962
tri 1521 937 1541 957 ne
rect 1541 937 1640 957
tri 1541 928 1550 937 ne
rect 1550 928 1640 937
rect 1674 928 2344 962
rect 2378 957 2497 962
tri 2497 957 2505 965 nw
rect 2378 937 2477 957
tri 2477 937 2497 957 nw
rect 2378 928 2465 937
tri 1550 925 1553 928 ne
rect 1553 925 2465 928
tri 2465 925 2477 937 nw
tri 4842 925 4854 937 se
rect 4854 925 4900 937
tri 1553 922 1556 925 ne
rect 1556 922 2462 925
tri 2462 922 2465 925 nw
tri 4839 922 4842 925 se
rect 4842 922 4860 925
tri 1556 908 1570 922 ne
rect 1570 908 2448 922
tri 2448 908 2462 922 nw
tri 2599 908 2613 922 se
rect 2613 916 4860 922
rect 2613 908 3984 916
rect 679 896 810 908
rect 679 862 685 896
rect 719 862 810 896
tri 1570 891 1587 908 ne
rect 1587 891 2431 908
tri 2431 891 2448 908 nw
tri 2582 891 2599 908 se
rect 2599 891 3984 908
tri 1587 890 1588 891 ne
rect 1588 890 2404 891
tri 1588 864 1614 890 ne
rect 1614 864 1640 890
rect 679 824 810 862
tri 1614 856 1622 864 ne
rect 1622 856 1640 864
rect 1674 856 2344 890
rect 2378 864 2404 890
tri 2404 864 2431 891 nw
tri 2555 864 2582 891 se
rect 2582 879 3984 891
rect 2582 864 2613 879
tri 2613 864 2628 879 nw
tri 3950 864 3965 879 ne
rect 3965 864 3984 879
rect 4036 891 4860 916
rect 4894 891 4900 925
rect 4036 879 4900 891
rect 4036 864 4055 879
tri 4055 864 4070 879 nw
tri 4820 864 4835 879 ne
rect 4835 864 4900 879
rect 2378 856 2393 864
tri 1622 853 1625 856 ne
rect 1625 853 2393 856
tri 2393 853 2404 864 nw
tri 2544 853 2555 864 se
rect 2555 853 2602 864
tri 2602 853 2613 864 nw
tri 3965 853 3976 864 ne
rect 3976 853 4044 864
tri 4044 853 4055 864 nw
tri 4835 853 4846 864 ne
rect 4846 853 4900 864
tri 1625 844 1634 853 ne
rect 1634 844 2384 853
tri 2384 844 2393 853 nw
tri 2535 844 2544 853 se
rect 2544 844 2588 853
tri 2530 839 2535 844 se
rect 2535 839 2588 844
tri 2588 839 2602 853 nw
tri 3976 851 3978 853 ne
rect 3978 852 4036 853
rect 3978 851 3984 852
tri 2528 837 2530 839 se
rect 2530 837 2586 839
tri 2586 837 2588 839 nw
tri 2521 830 2528 837 se
rect 2528 830 2579 837
tri 2579 830 2586 837 nw
rect 2987 830 3033 842
rect 679 790 685 824
rect 719 790 810 824
tri 2500 809 2521 830 se
rect 2521 809 2558 830
tri 2558 809 2579 830 nw
tri 2497 806 2500 809 se
rect 2500 806 2555 809
tri 2555 806 2558 809 nw
tri 2488 797 2497 806 se
rect 2497 797 2545 806
rect 679 778 810 790
rect 24 763 70 765
rect 21 757 73 763
rect 21 693 73 705
rect 1719 742 1771 748
rect 1841 745 1847 797
rect 1899 745 1911 797
rect 1963 791 2111 797
tri 2487 796 2488 797 se
rect 2488 796 2545 797
tri 2545 796 2555 806 nw
rect 2987 796 2993 830
rect 3027 796 3033 830
rect 1963 757 1993 791
rect 2027 757 2065 791
rect 2099 757 2111 791
tri 2474 783 2487 796 se
rect 2487 783 2532 796
tri 2532 783 2545 796 nw
rect 1963 751 2111 757
rect 2344 776 2525 783
tri 2525 776 2532 783 nw
rect 2344 767 2516 776
tri 2516 767 2525 776 nw
rect 2344 765 2514 767
tri 2514 765 2516 767 nw
rect 2344 758 2507 765
tri 2507 758 2514 765 nw
rect 2987 758 3033 796
rect 2344 751 2500 758
tri 2500 751 2507 758 nw
rect 1963 745 1975 751
tri 1975 745 1981 751 nw
rect 2344 748 2497 751
tri 2497 748 2500 751 nw
rect 2344 741 2490 748
tri 2490 741 2497 748 nw
rect 21 635 73 641
rect 326 689 372 701
tri 372 689 384 701 sw
tri 571 689 583 701 se
rect 583 689 629 701
tri 629 689 641 701 sw
tri 765 689 777 701 se
rect 777 689 823 701
rect 326 655 332 689
rect 366 674 384 689
tri 384 674 399 689 sw
tri 556 674 571 689 se
rect 571 674 589 689
rect 366 655 589 674
rect 623 674 641 689
tri 641 674 656 689 sw
tri 750 674 765 689 se
rect 765 674 783 689
rect 623 655 783 674
rect 817 655 823 689
rect 326 617 823 655
rect 326 583 332 617
rect 366 610 589 617
rect 366 583 379 610
tri 379 583 406 610 nw
tri 549 583 576 610 ne
rect 576 583 589 610
rect 623 610 783 617
rect 623 583 636 610
tri 636 583 663 610 nw
tri 744 583 771 610 ne
rect 771 583 783 610
rect 817 583 823 617
rect 1069 688 1347 697
tri 1347 688 1356 697 sw
rect 2987 724 2993 758
rect 3027 724 3033 758
rect 2987 712 3033 724
rect 3255 839 3301 842
tri 3301 839 3304 842 sw
rect 3255 837 3304 839
tri 3304 837 3306 839 sw
rect 3639 837 3685 849
rect 3255 834 3306 837
tri 3306 834 3309 837 sw
rect 3255 830 3309 834
rect 3255 796 3261 830
rect 3295 822 3309 830
tri 3309 822 3321 834 sw
tri 3627 822 3639 834 se
rect 3639 822 3645 837
rect 3295 809 3321 822
tri 3321 809 3334 822 sw
tri 3614 809 3627 822 se
rect 3627 809 3645 822
rect 3295 806 3334 809
tri 3334 806 3337 809 sw
tri 3611 806 3614 809 se
rect 3614 806 3645 809
rect 3295 803 3337 806
tri 3337 803 3340 806 sw
tri 3608 803 3611 806 se
rect 3611 803 3645 806
rect 3679 803 3685 837
rect 3295 802 3340 803
tri 3340 802 3341 803 sw
tri 3607 802 3608 803 se
rect 3608 802 3685 803
rect 3295 801 3341 802
tri 3341 801 3342 802 sw
tri 3606 801 3607 802 se
rect 3607 801 3685 802
rect 3295 800 3342 801
tri 3342 800 3343 801 sw
tri 3605 800 3606 801 se
rect 3606 800 3685 801
rect 3295 796 3685 800
rect 3255 765 3685 796
rect 3255 758 3645 765
rect 3255 724 3261 758
rect 3295 754 3645 758
rect 3295 751 3332 754
tri 3332 751 3335 754 nw
tri 3605 751 3608 754 ne
rect 3608 751 3645 754
rect 3295 748 3329 751
tri 3329 748 3332 751 nw
tri 3608 748 3611 751 ne
rect 3611 748 3645 751
rect 3295 741 3322 748
tri 3322 741 3329 748 nw
tri 3611 741 3618 748 ne
rect 3618 741 3645 748
rect 3295 731 3312 741
tri 3312 731 3322 741 nw
tri 3618 731 3628 741 ne
rect 3628 731 3645 741
rect 3679 731 3685 765
rect 3295 724 3302 731
rect 3255 721 3302 724
tri 3302 721 3312 731 nw
tri 3628 721 3638 731 ne
rect 3638 721 3685 731
rect 3731 839 3777 851
tri 3978 845 3984 851 ne
rect 3731 805 3737 839
rect 3771 805 3777 839
rect 3731 783 3777 805
tri 3777 783 3795 801 sw
tri 4036 845 4044 853 nw
tri 4846 851 4848 853 ne
rect 4848 851 4860 853
rect 4115 839 4161 851
tri 4848 845 4854 851 ne
rect 4115 805 4121 839
rect 4155 805 4161 839
rect 4854 819 4860 851
rect 4894 819 4900 853
rect 5751 829 5918 985
rect 4854 807 4900 819
rect 4937 812 4989 822
rect 3984 794 4036 800
tri 4108 794 4115 801 se
rect 4115 794 4161 805
tri 4097 783 4108 794 se
rect 4108 783 4161 794
tri 4918 783 4937 802 se
rect 3731 781 3795 783
tri 3795 781 3797 783 sw
tri 4095 781 4097 783 se
rect 4097 781 4161 783
tri 4916 781 4918 783 se
rect 4918 781 4937 783
rect 3731 776 3797 781
tri 3797 776 3802 781 sw
tri 4090 776 4095 781 se
rect 4095 776 4161 781
rect 3731 767 3802 776
tri 3802 767 3811 776 sw
tri 4081 767 4090 776 se
rect 4090 767 4161 776
rect 3731 733 3737 767
rect 3771 766 3811 767
tri 3811 766 3812 767 sw
tri 4080 766 4081 767 se
rect 4081 766 4121 767
rect 3771 733 4121 766
rect 4155 733 4161 767
rect 3731 721 4161 733
rect 4210 776 4675 781
tri 4675 776 4680 781 sw
tri 4911 776 4916 781 se
rect 4916 776 4937 781
rect 4210 760 4937 776
tri 7318 767 7360 809 ne
rect 4210 748 4989 760
rect 4210 747 4937 748
rect 4210 741 4272 747
tri 4272 741 4278 747 nw
tri 4619 742 4624 747 ne
rect 4624 742 4937 747
tri 4909 741 4910 742 ne
rect 4910 741 4937 742
rect 4210 738 4269 741
tri 4269 738 4272 741 nw
tri 4910 738 4913 741 ne
rect 4913 738 4937 741
rect 4210 725 4256 738
tri 4256 725 4269 738 nw
tri 4913 725 4926 738 ne
rect 4926 725 4937 738
tri 4206 721 4210 725 se
rect 4210 721 4245 725
rect 3255 712 3301 721
tri 3301 720 3302 721 nw
tri 3638 720 3639 721 ne
rect 3639 719 3685 721
tri 4204 719 4206 721 se
rect 4206 719 4245 721
tri 4200 715 4204 719 se
rect 4204 715 4245 719
rect 1719 688 1728 690
rect 1762 688 1771 690
rect 1069 685 1356 688
rect 1069 651 1075 685
rect 1109 663 1356 685
tri 1356 663 1381 688 sw
rect 1719 678 1771 688
rect 1109 651 1381 663
rect 1069 650 1381 651
tri 1381 650 1394 663 sw
rect 1069 616 1394 650
tri 1394 616 1428 650 sw
rect 1719 616 1728 626
rect 1762 616 1771 626
rect 1069 613 1428 616
rect 326 579 375 583
tri 375 579 379 583 nw
tri 576 579 580 583 ne
rect 580 579 632 583
tri 632 579 636 583 nw
tri 771 579 775 583 ne
rect 775 579 823 583
rect 326 571 372 579
tri 372 576 375 579 nw
tri 580 576 583 579 ne
rect 583 571 629 579
tri 629 576 632 579 nw
tri 775 577 777 579 ne
rect 777 571 823 579
rect 980 574 1026 586
rect -65 539 -13 545
rect -65 473 -13 487
rect -65 415 -13 421
rect 110 539 162 545
rect 980 540 986 574
rect 1020 540 1026 574
rect 1069 579 1075 613
rect 1109 607 1428 613
tri 1428 607 1437 616 sw
rect 1109 604 1437 607
tri 1437 604 1440 607 sw
rect 1719 604 1771 616
rect 2887 707 2933 709
tri 2933 707 2935 709 sw
tri 3079 707 3081 709 se
rect 3081 707 3127 709
tri 3127 707 3129 709 sw
tri 3337 707 3339 709 se
rect 3339 707 3385 709
rect 2887 697 2935 707
tri 2935 697 2945 707 sw
tri 3069 697 3079 707 se
rect 3079 697 3129 707
tri 3129 697 3139 707 sw
tri 3327 697 3337 707 se
rect 3337 697 3385 707
rect 2887 663 2893 697
rect 2927 682 2945 697
tri 2945 682 2960 697 sw
tri 3054 682 3069 697 se
rect 3069 682 3087 697
rect 2927 663 3087 682
rect 3121 682 3139 697
tri 3139 682 3154 697 sw
tri 3312 682 3327 697 se
rect 3327 682 3345 697
rect 3121 663 3345 682
rect 3379 663 3385 697
rect 3474 663 3480 715
rect 3532 663 3544 715
rect 3596 714 3602 715
tri 3602 714 3603 715 sw
tri 4199 714 4200 715 se
rect 4200 714 4245 715
tri 4245 714 4256 725 nw
tri 4926 719 4932 725 ne
rect 4932 719 4937 725
rect 3596 707 3603 714
tri 3603 707 3610 714 sw
tri 4192 707 4199 714 se
rect 4199 707 4244 714
tri 4244 713 4245 714 nw
rect 3596 691 3610 707
tri 3610 691 3626 707 sw
tri 4176 691 4192 707 se
rect 4192 691 4244 707
rect 3596 663 4244 691
rect 4468 707 4514 719
tri 4932 714 4937 719 ne
rect 4468 673 4474 707
rect 4508 673 4514 707
rect 7360 714 7412 809
tri 7412 767 7454 809 nw
rect 4937 690 4989 696
tri 4462 663 4468 669 se
rect 4468 663 4514 673
rect 2887 625 3385 663
tri 4434 635 4462 663 se
rect 4462 635 4514 663
rect 1109 591 1440 604
tri 1440 591 1453 604 sw
rect 2887 591 2893 625
rect 2927 618 3087 625
rect 2927 604 2953 618
tri 2953 604 2967 618 nw
tri 3047 604 3061 618 ne
rect 3061 604 3087 618
rect 2927 591 2940 604
tri 2940 591 2953 604 nw
tri 3061 591 3074 604 ne
rect 3074 591 3087 604
rect 3121 618 3345 625
rect 3121 591 3134 618
tri 3134 591 3161 618 nw
tri 3305 591 3332 618 ne
rect 3332 591 3345 618
rect 3379 591 3385 625
rect 1109 579 1453 591
rect 1069 567 1453 579
tri 1453 567 1477 591 sw
rect 2887 579 2933 591
tri 2933 584 2940 591 nw
tri 3074 584 3081 591 ne
rect 3081 579 3127 591
tri 3127 584 3134 591 nw
tri 3332 584 3339 591 ne
rect 3339 579 3385 591
rect 3425 601 4474 635
rect 4508 601 4514 635
rect 3425 574 3466 601
tri 3466 574 3493 601 nw
tri 4456 589 4468 601 ne
rect 4468 589 4514 601
tri 1293 562 1298 567 ne
rect 1298 562 1477 567
tri 1477 562 1482 567 sw
tri 1298 559 1301 562 ne
rect 1301 559 1482 562
tri 1482 559 1485 562 sw
tri 1301 555 1305 559 ne
rect 1305 555 1485 559
tri 1485 555 1489 559 sw
tri 1305 553 1307 555 ne
rect 1307 553 1489 555
tri 1489 553 1491 555 sw
rect 110 473 162 487
rect 110 415 162 421
rect 415 526 461 538
rect 415 492 421 526
rect 455 521 461 526
tri 461 521 478 538 sw
tri 963 521 980 538 se
rect 980 521 1026 540
tri 1307 521 1339 553 ne
rect 1339 547 1520 553
rect 1339 521 1468 547
rect 455 504 478 521
tri 478 504 495 521 sw
tri 946 504 963 521 se
rect 963 504 1026 521
rect 455 502 1026 504
rect 455 492 986 502
rect 415 470 986 492
rect 415 468 489 470
tri 489 468 491 470 nw
tri 966 468 968 470 ne
rect 968 468 986 470
rect 1020 468 1026 502
tri 1339 490 1370 521 ne
rect 1370 495 1468 521
tri 3400 521 3425 546 se
rect 3425 521 3459 574
tri 3459 567 3466 574 nw
tri 3391 512 3400 521 se
rect 3400 512 3459 521
rect 1370 490 1520 495
tri 1370 487 1373 490 ne
rect 1373 487 1520 490
tri 1373 483 1377 487 ne
rect 1377 483 1520 487
rect 415 456 477 468
tri 477 456 489 468 nw
tri 968 456 980 468 ne
rect 980 456 1026 468
tri 1377 456 1404 483 ne
rect 1404 481 1520 483
rect 1404 456 1468 481
rect 415 455 476 456
tri 476 455 477 456 nw
tri 1404 455 1405 456 ne
rect 1405 455 1468 456
rect 415 454 461 455
rect 415 420 421 454
rect 455 420 461 454
tri 461 440 476 455 nw
tri 1405 440 1420 455 ne
rect 1420 440 1468 455
tri 1420 423 1437 440 ne
rect 1437 429 1468 440
rect 1437 423 1520 429
rect 1840 455 2566 461
rect 3257 460 3263 512
rect 3315 460 3327 512
rect 3379 460 3459 512
rect 3550 561 3602 567
rect 3550 494 3602 509
rect 415 408 461 420
rect 1840 421 1852 455
rect 1886 421 1924 455
rect 1958 421 2448 455
rect 2482 421 2520 455
rect 2554 421 2566 455
rect 3550 436 3602 442
rect 4027 561 4079 567
rect 4027 494 4079 509
rect 4027 436 4079 442
rect 4200 561 4252 567
rect 4200 494 4252 509
rect 4200 436 4252 442
rect 4383 565 4435 571
rect 4383 498 4435 513
rect 4383 440 4435 446
rect 4552 565 4604 571
rect 4552 498 4604 513
rect 5024 568 5076 574
rect 5024 504 5076 516
rect 5024 446 5076 452
rect 4552 440 4604 446
rect 5027 444 5073 446
rect 1840 415 2566 421
rect 1452 378 2178 384
rect 1452 344 1464 378
rect 1498 344 1536 378
rect 1570 344 2060 378
rect 2094 344 2132 378
rect 2166 344 2178 378
rect 1452 338 2178 344
tri 2777 338 2785 346 se
rect 2785 345 5202 346
rect 2785 338 3730 345
tri 2776 337 2777 338 se
rect 2777 337 3730 338
rect -185 333 1250 337
tri 1250 333 1254 337 sw
tri 2772 333 2776 337 se
rect 2776 333 3730 337
rect -185 325 1254 333
rect -185 291 210 325
rect 244 291 510 325
rect 544 291 862 325
rect 896 291 1162 325
rect 1196 310 1254 325
tri 1254 310 1277 333 sw
tri 2761 322 2772 333 se
rect 2772 322 2817 333
tri 2488 316 2494 322 se
rect 2494 316 2518 322
rect 2211 310 2518 316
rect 1196 306 1277 310
tri 1277 306 1281 310 sw
rect 1196 291 1634 306
rect -185 261 1634 291
rect 2211 276 2223 310
rect 2257 276 2295 310
rect 2329 276 2518 310
tri 1634 261 1644 271 sw
rect 2211 270 2518 276
rect 2570 270 2582 322
rect 2634 270 2640 322
tri 2738 299 2761 322 se
rect 2761 299 2817 322
rect 2851 299 3169 333
rect 3203 299 3469 333
rect 3503 299 3730 333
tri 2709 270 2738 299 se
rect 2738 293 3730 299
rect 3782 293 3808 345
rect 3860 293 3887 345
rect 3939 333 5202 345
rect 3939 299 4297 333
rect 4331 299 4773 333
rect 4807 299 5202 333
rect 3939 293 5202 299
rect 2738 270 5202 293
tri 2700 261 2709 270 se
rect 2709 266 5202 270
rect 2709 261 3730 266
rect -185 253 1644 261
rect -185 219 210 253
rect 244 219 510 253
rect 544 219 862 253
rect 896 219 1162 253
rect 1196 242 1644 253
tri 1644 242 1663 261 sw
tri 2681 242 2700 261 se
rect 2700 242 2817 261
rect 1196 230 2817 242
rect 1196 219 1640 230
rect -185 196 1640 219
rect 1674 196 2344 230
rect 2378 227 2817 230
rect 2851 227 3169 261
rect 3203 227 3469 261
rect 3503 227 3730 261
rect 2378 214 3730 227
rect 3782 214 3808 266
rect 3860 214 3887 266
rect 3939 261 5202 266
rect 3939 227 4297 261
rect 4331 227 4773 261
rect 4807 227 5202 261
rect 3939 214 5202 227
rect 2378 196 5202 214
rect -185 187 5202 196
rect -185 176 3730 187
rect 3782 176 3808 187
rect -185 158 2817 176
rect -185 151 1640 158
rect -185 122 337 151
tri 300 117 305 122 ne
rect 305 117 337 122
rect 371 117 409 151
rect 443 117 481 151
rect 515 117 553 151
rect 587 117 625 151
rect 659 117 697 151
rect 731 117 769 151
rect 803 117 841 151
rect 875 117 913 151
rect 947 117 985 151
rect 1019 117 1057 151
rect 1091 117 1129 151
rect 1163 117 1201 151
rect 1235 124 1640 151
rect 1674 124 2344 158
rect 2378 142 2817 158
rect 2851 142 2889 176
rect 2923 142 2961 176
rect 2995 142 3033 176
rect 3067 142 3105 176
rect 3139 142 3177 176
rect 3211 142 3249 176
rect 3283 142 3321 176
rect 3355 142 3393 176
rect 3427 142 3465 176
rect 3499 142 3537 176
rect 3571 142 3609 176
rect 3643 142 3681 176
rect 3715 142 3730 176
rect 3787 142 3808 176
rect 2378 135 3730 142
rect 3782 135 3808 142
rect 3860 135 3887 187
rect 3939 176 5202 187
rect 3939 142 3969 176
rect 4003 142 4041 176
rect 4075 142 4113 176
rect 4147 142 4185 176
rect 4219 142 4257 176
rect 4291 142 4329 176
rect 4363 142 4401 176
rect 4435 142 4473 176
rect 4507 142 4545 176
rect 4579 142 4617 176
rect 4651 142 4689 176
rect 4723 142 4761 176
rect 4795 142 4833 176
rect 4867 142 4905 176
rect 4939 142 4977 176
rect 5011 142 5049 176
rect 5083 142 5121 176
rect 5155 142 5202 176
rect 3939 135 5202 142
rect 2378 130 5202 135
rect 2378 124 2805 130
rect 1235 117 2805 124
tri 305 105 317 117 ne
rect 317 112 2805 117
tri 2805 112 2823 130 nw
rect 317 105 1247 112
tri 1247 105 1254 112 nw
<< via1 >>
rect 2706 2797 2758 2849
rect 2777 2797 2829 2849
rect 3932 2797 3984 2849
rect 3996 2797 4048 2849
rect 31 2705 83 2757
rect 95 2705 147 2757
rect 2486 2705 2538 2757
rect 2550 2705 2602 2757
rect 129 2613 181 2665
rect 193 2613 245 2665
rect 2064 2613 2116 2665
rect 2128 2613 2180 2665
rect 3443 2613 3495 2665
rect 3507 2613 3559 2665
rect 4482 2613 4534 2665
rect 4546 2613 4598 2665
rect -133 2521 -81 2573
rect -69 2521 -17 2573
rect 1681 2521 1733 2573
rect 1745 2521 1797 2573
rect 4313 2521 4365 2573
rect 4377 2521 4429 2573
rect 1413 2429 1465 2481
rect 1477 2429 1529 2481
rect 4867 2429 4919 2481
rect 4931 2429 4983 2481
rect 1873 2337 1925 2389
rect 1937 2337 1989 2389
rect 4221 2337 4273 2389
rect 4285 2337 4337 2389
rect -63 1850 -11 1856
rect -63 1816 -54 1850
rect -54 1816 -20 1850
rect -20 1816 -11 1850
rect -63 1804 -11 1816
rect -63 1778 -11 1792
rect -63 1744 -54 1778
rect -54 1744 -20 1778
rect -20 1744 -11 1778
rect -63 1740 -11 1744
rect 123 1850 175 1856
rect 123 1816 132 1850
rect 132 1816 166 1850
rect 166 1816 175 1850
rect 123 1804 175 1816
rect 123 1778 175 1792
rect 123 1744 132 1778
rect 132 1744 166 1778
rect 166 1744 175 1778
rect 123 1740 175 1744
rect 1585 1781 1637 1833
rect 1585 1717 1637 1769
rect 3257 1842 3309 1848
rect 3257 1808 3267 1842
rect 3267 1808 3301 1842
rect 3301 1808 3309 1842
rect 3257 1796 3309 1808
rect 3257 1770 3309 1777
rect 2048 1712 2100 1764
rect 2112 1712 2164 1764
rect 2524 1695 2576 1747
rect 3257 1736 3267 1770
rect 3267 1736 3301 1770
rect 3301 1736 3309 1770
rect 3466 1829 3518 1881
rect 3466 1765 3518 1817
rect 3630 1846 3682 1898
rect 3630 1782 3682 1834
rect 4467 1833 4519 1885
rect 4467 1767 4519 1819
rect 3257 1725 3309 1736
rect 2524 1631 2576 1683
rect 4101 1682 4153 1734
rect 4165 1682 4217 1734
rect 3984 1643 4036 1649
rect 3984 1609 3997 1643
rect 3997 1609 4031 1643
rect 4031 1609 4036 1643
rect 3984 1597 4036 1609
rect 3984 1571 4036 1583
rect 3984 1537 3997 1571
rect 3997 1537 4031 1571
rect 4031 1537 4036 1571
rect 3984 1531 4036 1537
rect 4200 1582 4252 1634
rect 4200 1518 4252 1570
rect 201 1477 253 1483
rect 201 1443 210 1477
rect 210 1443 244 1477
rect 244 1443 253 1477
rect 201 1431 253 1443
rect 201 1405 253 1417
rect 201 1371 210 1405
rect 210 1371 244 1405
rect 244 1371 253 1405
rect 201 1365 253 1371
rect 410 1484 462 1493
rect 410 1450 421 1484
rect 421 1450 455 1484
rect 455 1450 462 1484
rect 410 1441 462 1450
rect 410 1412 462 1424
rect 410 1378 421 1412
rect 421 1378 455 1412
rect 455 1378 462 1412
rect 4291 1492 4343 1544
rect 4291 1428 4343 1480
rect 410 1372 462 1378
rect 3984 864 4036 916
rect 21 753 73 757
rect 21 719 30 753
rect 30 719 64 753
rect 64 719 73 753
rect 21 705 73 719
rect 1847 745 1899 797
rect 1911 745 1963 797
rect 1719 722 1771 742
rect 21 681 73 693
rect 21 647 30 681
rect 30 647 64 681
rect 64 647 73 681
rect 21 641 73 647
rect 1719 690 1728 722
rect 1728 690 1762 722
rect 1762 690 1771 722
rect 3984 800 4036 852
rect 4937 810 4989 812
rect 4937 776 4949 810
rect 4949 776 4983 810
rect 4983 776 4989 810
rect 4937 760 4989 776
rect 4937 738 4989 748
rect 1719 650 1771 678
rect 1719 626 1728 650
rect 1728 626 1762 650
rect 1762 626 1771 650
rect -65 533 -13 539
rect -65 499 -56 533
rect -56 499 -22 533
rect -22 499 -13 533
rect -65 487 -13 499
rect -65 461 -13 473
rect -65 427 -56 461
rect -56 427 -22 461
rect -22 427 -13 461
rect -65 421 -13 427
rect 110 533 162 539
rect 3480 663 3532 715
rect 3544 663 3596 715
rect 4937 704 4949 738
rect 4949 704 4983 738
rect 4983 704 4989 738
rect 4937 696 4989 704
rect 110 499 119 533
rect 119 499 153 533
rect 153 499 162 533
rect 110 487 162 499
rect 110 461 162 473
rect 110 427 119 461
rect 119 427 153 461
rect 153 427 162 461
rect 110 421 162 427
rect 1468 495 1520 547
rect 1468 429 1520 481
rect 3263 460 3315 512
rect 3327 460 3379 512
rect 3550 555 3602 561
rect 3550 521 3559 555
rect 3559 521 3593 555
rect 3593 521 3602 555
rect 3550 509 3602 521
rect 3550 483 3602 494
rect 3550 449 3559 483
rect 3559 449 3593 483
rect 3593 449 3602 483
rect 3550 442 3602 449
rect 4027 555 4079 561
rect 4027 521 4036 555
rect 4036 521 4070 555
rect 4070 521 4079 555
rect 4027 509 4079 521
rect 4027 483 4079 494
rect 4027 449 4036 483
rect 4036 449 4070 483
rect 4070 449 4079 483
rect 4027 442 4079 449
rect 4200 555 4252 561
rect 4200 521 4209 555
rect 4209 521 4243 555
rect 4243 521 4252 555
rect 4200 509 4252 521
rect 4200 483 4252 494
rect 4200 449 4209 483
rect 4209 449 4243 483
rect 4243 449 4252 483
rect 4200 442 4252 449
rect 4383 559 4435 565
rect 4383 525 4392 559
rect 4392 525 4426 559
rect 4426 525 4435 559
rect 4383 513 4435 525
rect 4383 487 4435 498
rect 4383 453 4392 487
rect 4392 453 4426 487
rect 4426 453 4435 487
rect 4383 446 4435 453
rect 4552 559 4604 565
rect 4552 525 4561 559
rect 4561 525 4595 559
rect 4595 525 4604 559
rect 4552 513 4604 525
rect 4552 487 4604 498
rect 4552 453 4561 487
rect 4561 453 4595 487
rect 4595 453 4604 487
rect 4552 446 4604 453
rect 5024 562 5076 568
rect 5024 528 5033 562
rect 5033 528 5067 562
rect 5067 528 5076 562
rect 5024 516 5076 528
rect 5024 490 5076 504
rect 5024 456 5033 490
rect 5033 456 5067 490
rect 5067 456 5076 490
rect 5024 452 5076 456
rect 2518 270 2570 322
rect 2582 270 2634 322
rect 3730 293 3782 345
rect 3808 293 3860 345
rect 3887 293 3939 345
rect 3730 214 3782 266
rect 3808 214 3860 266
rect 3887 214 3939 266
rect 3730 176 3782 187
rect 3808 176 3860 187
rect 3730 142 3753 176
rect 3753 142 3782 176
rect 3808 142 3825 176
rect 3825 142 3859 176
rect 3859 142 3860 176
rect 3730 135 3782 142
rect 3808 135 3860 142
rect 3887 176 3939 187
rect 3887 142 3897 176
rect 3897 142 3931 176
rect 3931 142 3939 176
rect 3887 135 3939 142
<< metal2 >>
tri 1744 2797 1796 2849 se
rect 1796 2797 2706 2849
rect 2758 2797 2777 2849
rect 2829 2797 2835 2849
rect 3926 2797 3932 2849
rect 3984 2797 3996 2849
rect 4048 2797 4054 2849
tri 1722 2775 1744 2797 se
rect 1744 2775 1796 2797
tri 1796 2775 1818 2797 nw
tri 3946 2775 3968 2797 ne
rect 3968 2775 4032 2797
tri 4032 2775 4054 2797 nw
tri 1710 2763 1722 2775 se
rect 1722 2763 1784 2775
tri 1784 2763 1796 2775 nw
tri 3968 2763 3980 2775 ne
tri 1704 2757 1710 2763 se
rect 1710 2757 1778 2763
tri 1778 2757 1784 2763 nw
rect 25 2705 31 2757
rect 83 2705 95 2757
rect 147 2705 153 2757
tri 1652 2705 1704 2757 se
rect 1704 2705 1726 2757
tri 1726 2705 1778 2757 nw
rect 2480 2705 2486 2757
rect 2538 2705 2550 2757
rect 2602 2705 2608 2757
rect 25 2701 107 2705
tri 107 2701 111 2705 nw
tri 1648 2701 1652 2705 se
rect 1652 2701 1722 2705
tri 1722 2701 1726 2705 nw
tri 2490 2701 2494 2705 ne
rect 2494 2701 2576 2705
rect -139 2521 -133 2573
rect -81 2521 -69 2573
rect -17 2521 -11 2573
tri -97 2487 -63 2521 ne
rect -63 1856 -11 2521
rect -63 1792 -11 1804
rect -63 1734 -11 1740
tri 9 1631 25 1647 se
rect 25 1631 77 2701
tri 77 2671 107 2701 nw
tri 1618 2671 1648 2701 se
rect 1648 2671 1686 2701
tri 1612 2665 1618 2671 se
rect 1618 2665 1686 2671
tri 1686 2665 1722 2701 nw
tri 2494 2671 2524 2701 ne
rect 123 2613 129 2665
rect 181 2613 193 2665
rect 245 2613 251 2665
tri 1585 2638 1612 2665 se
rect 1612 2638 1659 2665
tri 1659 2638 1686 2665 nw
rect 123 1856 175 2613
tri 175 2579 209 2613 nw
rect 1407 2429 1413 2481
rect 1465 2429 1477 2481
rect 1529 2429 1535 2481
tri 1434 2395 1468 2429 ne
rect 123 1792 175 1804
rect 123 1734 175 1740
tri 3 1625 9 1631 se
rect 9 1625 77 1631
tri -13 1609 3 1625 se
rect 3 1609 61 1625
tri 61 1609 77 1625 nw
tri -25 1597 -13 1609 se
rect -13 1597 49 1609
tri 49 1597 61 1609 nw
tri -39 1583 -25 1597 se
rect -25 1583 35 1597
tri 35 1583 49 1597 nw
tri -65 1557 -39 1583 se
rect -39 1557 -13 1583
rect -65 539 -13 1557
tri -13 1535 35 1583 nw
rect 410 1493 462 1499
rect 201 1483 253 1489
rect 201 1417 253 1431
rect 410 1424 462 1441
rect 410 1366 462 1372
tri 179 1154 201 1176 se
rect 201 1154 253 1365
tri 162 1137 179 1154 se
rect 179 1137 236 1154
tri 236 1137 253 1154 nw
tri 110 1085 162 1137 se
rect 21 757 73 763
rect 21 693 73 705
rect 21 635 73 641
rect -65 473 -13 487
rect -65 415 -13 421
rect 110 539 162 1085
tri 162 1063 236 1137 nw
rect 110 473 162 487
rect 1468 547 1520 2429
tri 1520 2414 1535 2429 nw
rect 1585 1833 1637 2638
tri 1637 2616 1659 2638 nw
rect 2058 2613 2064 2665
rect 2116 2613 2128 2665
rect 2180 2613 2186 2665
tri 2068 2579 2102 2613 ne
rect 1675 2521 1681 2573
rect 1733 2521 1745 2573
rect 1797 2521 1803 2573
tri 1685 2489 1717 2521 ne
rect 1717 2489 1771 2521
tri 1771 2489 1803 2521 nw
tri 1717 2487 1719 2489 ne
rect 1585 1769 1637 1781
rect 1585 1711 1637 1717
rect 1719 742 1771 2489
rect 1867 2337 1873 2389
rect 1925 2337 1937 2389
rect 1989 2337 1995 2389
tri 1867 2333 1871 2337 ne
tri 1844 800 1871 827 se
rect 1871 800 1917 2337
tri 1917 2303 1951 2337 nw
tri 2100 1796 2102 1798 se
rect 2102 1796 2148 2613
tri 2148 2581 2180 2613 nw
tri 2514 2429 2524 2439 se
rect 2524 2429 2576 2701
tri 2576 2673 2608 2705 nw
rect 3437 2613 3443 2665
rect 3495 2613 3507 2665
rect 3559 2613 3565 2665
tri 3437 2584 3466 2613 ne
tri 2490 2405 2514 2429 se
rect 2514 2405 2576 2429
rect 2434 2353 2576 2405
rect 2434 2337 2504 2353
tri 2504 2337 2520 2353 nw
rect 2434 2179 2486 2337
tri 2486 2319 2504 2337 nw
tri 2486 2179 2520 2213 sw
rect 2434 2127 2576 2179
tri 2490 2093 2524 2127 ne
tri 2081 1777 2100 1796 se
rect 2100 1777 2148 1796
tri 2148 1777 2157 1786 sw
tri 2068 1764 2081 1777 se
rect 2081 1764 2157 1777
tri 2157 1764 2170 1777 sw
rect 2042 1712 2048 1764
rect 2100 1712 2112 1764
rect 2164 1712 2170 1764
rect 2524 1747 2576 2127
rect 3466 1881 3518 2613
tri 3518 2579 3552 2613 nw
rect 3980 2521 4032 2775
rect 4476 2613 4482 2665
rect 4534 2613 4546 2665
rect 4598 2613 4604 2665
tri 4518 2579 4552 2613 ne
tri 4032 2521 4036 2525 sw
rect 4307 2521 4313 2573
rect 4365 2521 4377 2573
rect 4429 2521 4435 2573
rect 3980 2491 4036 2521
tri 4036 2491 4066 2521 sw
tri 4349 2491 4379 2521 ne
rect 4379 2491 4435 2521
rect 3980 2439 4143 2491
tri 4379 2487 4383 2491 ne
tri 4057 2429 4067 2439 ne
rect 4067 2429 4143 2439
tri 4067 2405 4091 2429 ne
rect 2524 1683 2576 1695
tri 1917 800 1948 831 sw
tri 1841 797 1844 800 se
rect 1844 797 1948 800
tri 1948 797 1951 800 sw
rect 1841 745 1847 797
rect 1899 745 1911 797
rect 1963 745 1969 797
rect 1719 678 1771 690
rect 1719 620 1771 626
rect 1468 481 1520 495
rect 1468 423 1520 429
rect 110 415 162 421
rect 2524 345 2576 1631
rect 3257 1848 3309 1854
rect 3257 1777 3309 1796
rect 3466 1817 3518 1829
rect 3466 1759 3518 1765
rect 3630 1898 3682 1904
rect 3630 1834 3682 1846
rect 3257 512 3309 1725
rect 3474 663 3480 715
rect 3532 663 3544 715
rect 3596 663 3602 715
tri 3562 568 3630 636 se
rect 3630 568 3682 1782
rect 4091 1767 4143 2429
rect 4215 2337 4221 2389
rect 4273 2337 4285 2389
rect 4337 2337 4343 2389
tri 4257 2303 4291 2337 ne
tri 4143 1767 4144 1768 sw
rect 4091 1734 4144 1767
tri 4144 1734 4177 1767 sw
rect 4091 1682 4101 1734
rect 4153 1682 4165 1734
rect 4217 1682 4223 1734
rect 3984 1649 4036 1655
rect 3984 1583 4036 1597
rect 3984 916 4036 1531
rect 3984 852 4036 864
rect 3984 794 4036 800
tri 3561 567 3562 568 se
rect 3562 567 3682 568
rect 3550 561 3682 567
tri 3309 512 3343 546 sw
rect 3257 460 3263 512
rect 3315 460 3327 512
rect 3379 460 3385 512
rect 3602 528 3682 561
tri 4027 614 4091 678 se
rect 4091 656 4143 1682
tri 4143 1648 4177 1682 nw
rect 4091 614 4101 656
tri 4101 614 4143 656 nw
rect 4200 1634 4252 1640
rect 4200 1570 4252 1582
rect 4027 561 4079 614
tri 4079 592 4101 614 nw
rect 3602 509 3639 528
tri 3639 509 3658 528 nw
rect 3550 504 3634 509
tri 3634 504 3639 509 nw
rect 3550 498 3628 504
tri 3628 498 3634 504 nw
rect 3550 494 3624 498
tri 3624 494 3628 498 nw
rect 4027 494 4079 509
tri 3602 472 3624 494 nw
tri 2576 345 2587 356 sw
tri 2512 322 2524 334 se
rect 2524 322 2587 345
tri 2587 322 2610 345 sw
rect 2512 270 2518 322
rect 2570 270 2582 322
rect 2634 270 2640 322
rect 3550 285 3602 442
rect 3724 345 3945 346
rect 3724 293 3730 345
rect 3782 293 3808 345
rect 3860 293 3887 345
rect 3939 293 3945 345
rect 3724 266 3945 293
rect 4027 269 4079 442
rect 4200 561 4252 1518
rect 4291 1544 4343 2337
rect 4291 1480 4343 1492
rect 4291 1422 4343 1428
rect 4200 494 4252 509
rect 4200 285 4252 442
rect 4383 565 4435 2491
rect 4383 498 4435 513
rect 4383 440 4435 446
rect 4467 1885 4519 1891
rect 4467 1819 4519 1833
rect 4467 305 4519 1767
rect 4552 565 4604 2613
rect 4861 2429 4867 2481
rect 4919 2429 4931 2481
rect 4983 2429 4989 2481
tri 4903 2395 4937 2429 ne
rect 4937 812 4989 2429
rect 4937 748 4989 760
rect 4937 690 4989 696
rect 4552 498 4604 513
rect 4552 440 4604 446
rect 5024 568 5076 587
rect 5024 504 5076 516
rect 5024 412 5076 452
rect 3724 214 3730 266
rect 3782 214 3808 266
rect 3860 214 3887 266
rect 3939 214 3945 266
rect 3724 187 3945 214
rect 3724 135 3730 187
rect 3782 135 3808 187
rect 3860 135 3887 187
rect 3939 135 3945 187
rect 3724 134 3945 135
use sky130_fd_io__com_ctl_ls_octl  sky130_fd_io__com_ctl_ls_octl_0
timestamp 1686671242
transform 1 0 5445 0 -1 2130
box -71 10 2077 2019
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1686671242
transform 1 0 3095 0 -1 2174
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1686671242
transform 1 0 3095 0 1 106
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_2
timestamp 1686671242
transform -1 0 618 0 1 98
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_3
timestamp 1686671242
transform -1 0 1270 0 1 98
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_4
timestamp 1686671242
transform -1 0 618 0 -1 2182
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1_i2c_fix  sky130_fd_io__hvsbt_inv_x1_i2c_fix_0
timestamp 1686671242
transform 1 0 2032 0 -1 3724
box 107 226 240 751
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_0
timestamp 1686671242
transform 1 0 2743 0 -1 2174
box 107 226 460 873
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_1
timestamp 1686671242
transform -1 0 3277 0 1 106
box 107 226 460 873
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_2
timestamp 1686671242
transform -1 0 970 0 -1 2182
box 107 226 460 873
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_3
timestamp 1686671242
transform -1 0 970 0 1 98
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1686671242
transform 1 0 3747 0 -1 2174
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1686671242
transform -1 0 3929 0 -1 2174
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_2
timestamp 1686671242
transform -1 0 4757 0 -1 2174
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_3
timestamp 1686671242
transform 1 0 4699 0 1 106
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_4
timestamp 1686671242
transform -1 0 4405 0 1 106
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_5
timestamp 1686671242
transform 1 0 3395 0 1 106
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_6
timestamp 1686671242
transform 1 0 4223 0 1 106
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_7
timestamp 1686671242
transform -1 0 318 0 1 98
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1686671242
transform 1 0 4699 0 -1 2174
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1686671242
transform 1 0 788 0 -1 2182
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_2
timestamp 1686671242
transform 1 0 -216 0 -1 2182
box 107 226 460 873
use sky130_fd_io__hvsbt_xor  sky130_fd_io__hvsbt_xor_0
timestamp 1686671242
transform -1 0 2723 0 1 -63
box 213 167 1215 838
use sky130_fd_io__hvsbt_xor  sky130_fd_io__hvsbt_xor_1
timestamp 1686671242
transform -1 0 2756 0 -1 2346
box 213 167 1215 838
<< labels >>
flabel metal2 s 27 664 64 728 3 FreeSans 520 0 0 0 PDEN_H_N[2]
port 2 nsew
flabel metal2 s 5032 478 5063 543 3 FreeSans 520 0 0 0 VREG_EN_H_N
port 1 nsew
flabel metal2 s 416 1379 454 1471 3 FreeSans 520 0 0 0 PUEN_0_H
port 3 nsew
flabel metal2 s 3554 290 3598 339 3 FreeSans 520 90 0 0 DM_H_N[0]
port 8 nsew
flabel metal2 s 4209 296 4244 341 3 FreeSans 520 90 0 0 DM_H_N[2]
port 10 nsew
flabel metal2 s 3989 891 4020 985 3 FreeSans 520 180 0 0 PUEN_2OR1_H
port 9 nsew
flabel metal2 s 4385 471 4434 524 3 FreeSans 520 90 0 0 DM_H[1]
port 4 nsew
flabel metal2 s 4553 463 4602 526 3 FreeSans 520 90 0 0 DM_H[0]
port 5 nsew
flabel metal2 s 2538 336 2564 385 3 FreeSans 520 90 0 0 DM_H[2]
port 6 nsew
flabel metal2 s 4036 297 4070 346 3 FreeSans 520 90 0 0 DM_H_N[1]
port 7 nsew
flabel metal2 s 3576 314 3576 314 3 FreeSans 520 90 0 0 DM_H_N[0]
flabel metal2 s 4004 938 4004 938 3 FreeSans 520 180 0 0 PUEN_2OR1_H
flabel metal2 s 4227 318 4227 318 3 FreeSans 520 90 0 0 DM_H_N[2]
flabel comment s 4058 183 4058 183 0 FreeSans 440 90 0 0 DM_H_N[1]
flabel comment s 4586 866 4586 866 0 FreeSans 440 270 0 0 DM_H[0]
flabel comment s 4408 849 4408 849 0 FreeSans 440 270 0 0 DM_H[1]
flabel comment s 5067 1248 5067 1248 0 FreeSans 440 90 0 0 DM_H[2]
flabel comment s 4234 179 4234 179 0 FreeSans 440 90 0 0 DM_H_N[2]
flabel comment s 3582 245 3582 245 0 FreeSans 440 270 0 0 DM_H_N[0]
flabel metal1 s 682 1761 722 1838 3 FreeSans 520 0 0 0 PUEN_H[0]
port 11 nsew
flabel metal1 s 5751 829 5918 985 3 FreeSans 520 180 0 0 VGND
port 18 nsew
flabel metal1 s 5540 1805 5851 2006 3 FreeSans 520 180 0 0 VCC_IO
port 14 nsew
flabel metal1 s 682 793 722 870 3 FreeSans 520 0 0 0 PUEN_H[1]
port 17 nsew
flabel metal1 s 7159 1677 7237 1745 3 FreeSans 520 0 0 0 VPWR
port 13 nsew
flabel metal1 s 5798 1449 5833 1488 3 FreeSans 520 0 0 0 SLOW_H
port 15 nsew
flabel metal1 s 6826 1452 6865 1496 3 FreeSans 520 0 0 0 HLD_I_H_N
port 12 nsew
flabel metal1 s 7159 1541 7237 1609 3 FreeSans 520 0 0 0 VPWR
port 13 nsew
flabel metal1 s 7371 1409 7459 1454 3 FreeSans 520 0 0 0 SLOW
port 20 nsew
flabel metal1 s 2192 3308 2231 3357 3 FreeSans 520 0 0 0 OD_H
port 19 nsew
flabel metal1 s 5483 1123 5522 1168 3 FreeSans 520 0 0 0 SLOW_H_N
port 16 nsew
flabel metal1 s 384 1005 695 1237 3 FreeSans 520 180 0 0 VCC_IO
port 14 nsew
flabel metal1 s 358 2015 525 2171 3 FreeSans 520 180 0 0 VGND
port 18 nsew
flabel metal1 s 2994 770 3024 830 3 FreeSans 520 180 0 0 PDEN_H_N[1]
port 21 nsew
flabel metal1 s 2992 1405 3026 1469 3 FreeSans 520 180 0 0 PDEN_H_N[0]
port 22 nsew
flabel metal1 s 2852 152 3019 322 3 FreeSans 520 180 0 0 VGND
port 18 nsew
flabel metal1 s 2851 1028 3162 1260 3 FreeSans 520 180 0 0 VCC_IO
port 14 nsew
flabel metal1 s 2852 2117 3019 2273 3 FreeSans 520 180 0 0 VGND
port 18 nsew
<< properties >>
string GDS_END 36671466
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 36598686
<< end >>
