magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 39 21 1011 203
rect 39 17 62 21
rect 28 -17 62 17
<< scnmos >>
rect 121 47 151 177
rect 200 47 230 177
rect 284 47 314 177
rect 368 47 398 177
rect 452 47 482 177
rect 524 47 554 177
rect 651 47 681 177
rect 735 47 765 177
rect 819 47 849 177
rect 903 47 933 177
<< scpmoshvt >>
rect 121 297 151 497
rect 200 297 230 497
rect 284 297 314 497
rect 368 297 398 497
rect 452 297 482 497
rect 524 297 554 497
rect 651 297 681 497
rect 735 297 765 497
rect 819 297 849 497
rect 903 297 933 497
<< ndiff >>
rect 65 161 121 177
rect 65 127 77 161
rect 111 127 121 161
rect 65 93 121 127
rect 65 59 77 93
rect 111 59 121 93
rect 65 47 121 59
rect 151 47 200 177
rect 230 93 284 177
rect 230 59 240 93
rect 274 59 284 93
rect 230 47 284 59
rect 314 47 368 177
rect 398 161 452 177
rect 398 127 408 161
rect 442 127 452 161
rect 398 93 452 127
rect 398 59 408 93
rect 442 59 452 93
rect 398 47 452 59
rect 482 47 524 177
rect 554 93 651 177
rect 554 59 588 93
rect 622 59 651 93
rect 554 47 651 59
rect 681 165 735 177
rect 681 131 691 165
rect 725 131 735 165
rect 681 97 735 131
rect 681 63 691 97
rect 725 63 735 97
rect 681 47 735 63
rect 765 93 819 177
rect 765 59 775 93
rect 809 59 819 93
rect 765 47 819 59
rect 849 165 903 177
rect 849 131 859 165
rect 893 131 903 165
rect 849 97 903 131
rect 849 63 859 97
rect 893 63 903 97
rect 849 47 903 63
rect 933 93 985 177
rect 933 59 943 93
rect 977 59 985 93
rect 933 47 985 59
<< pdiff >>
rect 47 477 121 497
rect 47 443 59 477
rect 93 443 121 477
rect 47 409 121 443
rect 47 375 59 409
rect 93 375 121 409
rect 47 341 121 375
rect 47 307 59 341
rect 93 307 121 341
rect 47 297 121 307
rect 151 297 200 497
rect 230 485 284 497
rect 230 451 240 485
rect 274 451 284 485
rect 230 297 284 451
rect 314 297 368 497
rect 398 411 452 497
rect 398 377 408 411
rect 442 377 452 411
rect 398 343 452 377
rect 398 309 408 343
rect 442 309 452 343
rect 398 297 452 309
rect 482 297 524 497
rect 554 485 651 497
rect 554 451 585 485
rect 619 451 651 485
rect 554 409 651 451
rect 554 375 585 409
rect 619 375 651 409
rect 554 341 651 375
rect 554 307 585 341
rect 619 307 651 341
rect 554 297 651 307
rect 681 485 735 497
rect 681 451 691 485
rect 725 451 735 485
rect 681 409 735 451
rect 681 375 691 409
rect 725 375 735 409
rect 681 341 735 375
rect 681 307 691 341
rect 725 307 735 341
rect 681 297 735 307
rect 765 485 819 497
rect 765 451 775 485
rect 809 451 819 485
rect 765 409 819 451
rect 765 375 775 409
rect 809 375 819 409
rect 765 297 819 375
rect 849 485 903 497
rect 849 451 859 485
rect 893 451 903 485
rect 849 409 903 451
rect 849 375 859 409
rect 893 375 903 409
rect 849 341 903 375
rect 849 307 859 341
rect 893 307 903 341
rect 849 297 903 307
rect 933 485 985 497
rect 933 451 943 485
rect 977 451 985 485
rect 933 409 985 451
rect 933 375 943 409
rect 977 375 985 409
rect 933 297 985 375
<< ndiffc >>
rect 77 127 111 161
rect 77 59 111 93
rect 240 59 274 93
rect 408 127 442 161
rect 408 59 442 93
rect 588 59 622 93
rect 691 131 725 165
rect 691 63 725 97
rect 775 59 809 93
rect 859 131 893 165
rect 859 63 893 97
rect 943 59 977 93
<< pdiffc >>
rect 59 443 93 477
rect 59 375 93 409
rect 59 307 93 341
rect 240 451 274 485
rect 408 377 442 411
rect 408 309 442 343
rect 585 451 619 485
rect 585 375 619 409
rect 585 307 619 341
rect 691 451 725 485
rect 691 375 725 409
rect 691 307 725 341
rect 775 451 809 485
rect 775 375 809 409
rect 859 451 893 485
rect 859 375 893 409
rect 859 307 893 341
rect 943 451 977 485
rect 943 375 977 409
<< poly >>
rect 121 497 151 523
rect 200 497 230 523
rect 284 497 314 523
rect 368 497 398 523
rect 452 497 482 523
rect 524 497 554 523
rect 651 497 681 523
rect 735 497 765 523
rect 819 497 849 523
rect 903 497 933 523
rect 121 265 151 297
rect 85 249 151 265
rect 85 215 101 249
rect 135 215 151 249
rect 85 199 151 215
rect 121 177 151 199
rect 200 265 230 297
rect 284 265 314 297
rect 200 249 314 265
rect 200 215 240 249
rect 274 215 314 249
rect 200 199 314 215
rect 200 177 230 199
rect 284 177 314 199
rect 368 265 398 297
rect 452 265 482 297
rect 368 249 482 265
rect 368 215 408 249
rect 442 215 482 249
rect 368 199 482 215
rect 368 177 398 199
rect 452 177 482 199
rect 524 265 554 297
rect 651 265 681 297
rect 735 265 765 297
rect 819 265 849 297
rect 903 265 933 297
rect 524 249 589 265
rect 524 215 539 249
rect 573 215 589 249
rect 524 199 589 215
rect 651 249 933 265
rect 651 215 691 249
rect 725 215 775 249
rect 809 215 859 249
rect 893 215 933 249
rect 651 199 933 215
rect 524 177 554 199
rect 651 177 681 199
rect 735 177 765 199
rect 819 177 849 199
rect 903 177 933 199
rect 121 21 151 47
rect 200 21 230 47
rect 284 21 314 47
rect 368 21 398 47
rect 452 21 482 47
rect 524 21 554 47
rect 651 21 681 47
rect 735 21 765 47
rect 819 21 849 47
rect 903 21 933 47
<< polycont >>
rect 101 215 135 249
rect 240 215 274 249
rect 408 215 442 249
rect 539 215 573 249
rect 691 215 725 249
rect 775 215 809 249
rect 859 215 893 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 477 93 493
rect 17 443 59 477
rect 224 485 290 527
rect 224 451 240 485
rect 274 451 290 485
rect 569 485 635 527
rect 17 409 93 443
rect 324 445 526 479
rect 324 417 358 445
rect 17 375 59 409
rect 17 341 93 375
rect 17 307 59 341
rect 17 291 93 307
rect 144 383 358 417
rect 17 177 51 291
rect 144 257 178 383
rect 392 377 408 411
rect 442 377 458 411
rect 392 349 458 377
rect 324 343 458 349
rect 85 249 178 257
rect 85 215 101 249
rect 135 215 178 249
rect 212 249 290 327
rect 212 215 240 249
rect 274 215 290 249
rect 324 309 408 343
rect 442 309 458 343
rect 324 177 358 309
rect 392 249 458 265
rect 392 215 408 249
rect 442 215 458 249
rect 492 249 526 445
rect 569 451 585 485
rect 619 451 635 485
rect 569 409 635 451
rect 569 375 585 409
rect 619 375 635 409
rect 569 341 635 375
rect 569 307 585 341
rect 619 307 635 341
rect 569 291 635 307
rect 675 485 741 493
rect 675 451 691 485
rect 725 451 741 485
rect 675 409 741 451
rect 675 375 691 409
rect 725 375 741 409
rect 675 341 741 375
rect 775 485 809 527
rect 775 409 809 451
rect 775 359 809 375
rect 843 485 909 493
rect 843 451 859 485
rect 893 451 909 485
rect 843 409 909 451
rect 843 375 859 409
rect 893 375 909 409
rect 675 307 691 341
rect 725 325 741 341
rect 843 341 909 375
rect 943 485 985 527
rect 977 451 985 485
rect 943 409 985 451
rect 977 375 985 409
rect 943 359 985 375
rect 843 325 859 341
rect 725 307 859 325
rect 893 325 909 341
rect 893 307 995 325
rect 675 291 995 307
rect 623 249 909 257
rect 492 215 539 249
rect 573 215 589 249
rect 623 215 691 249
rect 725 215 775 249
rect 809 215 859 249
rect 893 215 909 249
rect 623 177 657 215
rect 943 181 995 291
rect 17 161 657 177
rect 17 127 77 161
rect 111 132 408 161
rect 111 127 127 132
rect 17 93 127 127
rect 392 127 408 132
rect 442 143 657 161
rect 691 165 995 181
rect 442 127 458 143
rect 17 59 77 93
rect 111 59 127 93
rect 17 51 127 59
rect 224 93 290 98
rect 224 59 240 93
rect 274 59 290 93
rect 224 17 290 59
rect 392 93 458 127
rect 725 143 859 165
rect 725 131 741 143
rect 392 59 408 93
rect 442 59 458 93
rect 392 51 458 59
rect 572 93 641 109
rect 691 98 741 131
rect 843 131 859 143
rect 893 143 995 165
rect 893 131 909 143
rect 572 59 588 93
rect 622 59 641 93
rect 572 17 641 59
rect 675 97 741 98
rect 675 63 691 97
rect 725 63 741 97
rect 675 51 741 63
rect 775 93 809 109
rect 775 17 809 59
rect 843 97 909 131
rect 843 63 859 97
rect 893 63 909 97
rect 843 51 909 63
rect 943 93 977 109
rect 943 17 977 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel locali s 948 221 982 255 0 FreeSans 250 0 0 0 X
port 8 nsew signal output
flabel locali s 948 289 982 323 0 FreeSans 250 0 0 0 X
port 8 nsew signal output
flabel locali s 396 221 430 255 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 212 221 246 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 212 289 246 323 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 948 153 982 187 0 FreeSans 250 0 0 0 X
port 8 nsew signal output
flabel nwell s 28 527 62 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 28 -17 62 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 28 -17 62 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 28 527 62 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 maj3_4
rlabel metal1 s 0 -48 1012 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_END 1668080
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1660210
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 25.300 0.000 
<< end >>
