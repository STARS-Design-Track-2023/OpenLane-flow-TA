magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -66 449 3042 897
rect -66 377 1029 449
rect 1434 377 3042 449
<< pwell >>
rect 1089 313 1374 361
rect 4 217 426 241
rect 1089 217 2972 313
rect 4 43 2972 217
rect -26 -43 3002 43
<< mvnmos >>
rect 87 131 187 215
rect 243 131 343 215
rect 1168 251 1268 335
rect 542 107 642 191
rect 698 107 798 191
rect 858 107 958 191
rect 1000 107 1100 191
rect 1370 203 1470 287
rect 1545 137 1645 287
rect 1687 137 1787 287
rect 1889 203 1989 287
rect 2031 203 2131 287
rect 2173 203 2273 287
rect 2329 203 2429 287
rect 2610 203 2710 287
rect 2789 137 2889 287
<< mvpmos >>
rect 84 593 184 743
rect 240 593 340 743
rect 562 529 662 613
rect 718 529 818 613
rect 882 529 982 613
rect 1024 529 1124 613
rect 1218 529 1318 613
rect 1374 529 1474 613
rect 1553 515 1653 715
rect 1695 515 1795 715
rect 2352 659 2452 743
rect 1889 515 1989 599
rect 2031 515 2131 599
rect 2187 515 2287 599
rect 2618 519 2718 669
rect 2793 519 2893 719
<< mvndiff >>
rect 30 190 87 215
rect 30 156 42 190
rect 76 156 87 190
rect 30 131 87 156
rect 187 190 243 215
rect 187 156 198 190
rect 232 156 243 190
rect 187 131 243 156
rect 343 190 400 215
rect 1115 310 1168 335
rect 1115 276 1123 310
rect 1157 276 1168 310
rect 1115 251 1168 276
rect 1268 287 1348 335
rect 1268 251 1370 287
rect 343 156 354 190
rect 388 156 400 190
rect 343 131 400 156
rect 485 166 542 191
rect 485 132 497 166
rect 531 132 542 166
rect 485 107 542 132
rect 642 166 698 191
rect 642 132 653 166
rect 687 132 698 166
rect 642 107 698 132
rect 798 166 858 191
rect 798 132 813 166
rect 847 132 858 166
rect 798 107 858 132
rect 958 107 1000 191
rect 1100 155 1153 191
rect 1100 121 1111 155
rect 1145 121 1153 155
rect 1100 107 1153 121
rect 1290 203 1370 251
rect 1470 275 1545 287
rect 1470 241 1500 275
rect 1534 241 1545 275
rect 1470 203 1545 241
rect 1492 183 1545 203
rect 1492 149 1500 183
rect 1534 149 1545 183
rect 1492 137 1545 149
rect 1645 137 1687 287
rect 1787 275 1889 287
rect 1787 241 1821 275
rect 1855 241 1889 275
rect 1787 203 1889 241
rect 1989 203 2031 287
rect 2131 203 2173 287
rect 2273 262 2329 287
rect 2273 228 2284 262
rect 2318 228 2329 262
rect 2273 203 2329 228
rect 2429 262 2486 287
rect 2429 228 2440 262
rect 2474 228 2486 262
rect 2429 203 2486 228
rect 2553 262 2610 287
rect 2553 228 2565 262
rect 2599 228 2610 262
rect 2553 203 2610 228
rect 2710 279 2789 287
rect 2710 245 2744 279
rect 2778 245 2789 279
rect 2710 203 2789 245
rect 1787 137 1837 203
rect 2732 179 2789 203
rect 2732 145 2744 179
rect 2778 145 2789 179
rect 2732 137 2789 145
rect 2889 279 2946 287
rect 2889 245 2900 279
rect 2934 245 2946 279
rect 2889 179 2946 245
rect 2889 145 2900 179
rect 2934 145 2946 179
rect 2889 137 2946 145
<< mvpdiff >>
rect 31 731 84 743
rect 31 697 39 731
rect 73 697 84 731
rect 31 639 84 697
rect 31 605 39 639
rect 73 605 84 639
rect 31 593 84 605
rect 184 735 240 743
rect 184 701 195 735
rect 229 701 240 735
rect 184 635 240 701
rect 184 601 195 635
rect 229 601 240 635
rect 184 593 240 601
rect 340 731 393 743
rect 340 697 351 731
rect 385 697 393 731
rect 340 639 393 697
rect 340 605 351 639
rect 385 605 393 639
rect 1496 707 1553 715
rect 1496 673 1508 707
rect 1542 673 1553 707
rect 1496 638 1553 673
rect 1496 613 1508 638
rect 340 593 393 605
rect 455 588 562 613
rect 455 554 463 588
rect 497 554 562 588
rect 455 529 562 554
rect 662 588 718 613
rect 662 554 673 588
rect 707 554 718 588
rect 662 529 718 554
rect 818 588 882 613
rect 818 554 829 588
rect 863 554 882 588
rect 818 529 882 554
rect 982 529 1024 613
rect 1124 605 1218 613
rect 1124 571 1137 605
rect 1171 571 1218 605
rect 1124 529 1218 571
rect 1318 588 1374 613
rect 1318 554 1329 588
rect 1363 554 1374 588
rect 1318 529 1374 554
rect 1474 604 1508 613
rect 1542 604 1553 638
rect 1474 569 1553 604
rect 1474 535 1508 569
rect 1542 535 1553 569
rect 1474 529 1553 535
rect 1496 515 1553 529
rect 1653 515 1695 715
rect 1795 661 1867 715
rect 1795 627 1825 661
rect 1859 627 1867 661
rect 1795 599 1867 627
rect 2264 718 2352 743
rect 2264 684 2276 718
rect 2310 684 2352 718
rect 2264 659 2352 684
rect 2452 718 2505 743
rect 2452 684 2463 718
rect 2497 684 2505 718
rect 2740 707 2793 719
rect 2452 659 2505 684
rect 2740 673 2748 707
rect 2782 673 2793 707
rect 2740 669 2793 673
rect 2565 657 2618 669
rect 1795 515 1889 599
rect 1989 515 2031 599
rect 2131 579 2187 599
rect 2131 545 2142 579
rect 2176 545 2187 579
rect 2131 515 2187 545
rect 2287 577 2337 599
rect 2287 561 2344 577
rect 2287 527 2298 561
rect 2332 527 2344 561
rect 2287 515 2344 527
rect 2565 623 2573 657
rect 2607 623 2618 657
rect 2565 565 2618 623
rect 2565 531 2573 565
rect 2607 531 2618 565
rect 2565 519 2618 531
rect 2718 636 2793 669
rect 2718 602 2748 636
rect 2782 602 2793 636
rect 2718 565 2793 602
rect 2718 531 2748 565
rect 2782 531 2793 565
rect 2718 519 2793 531
rect 2893 707 2946 719
rect 2893 673 2904 707
rect 2938 673 2946 707
rect 2893 636 2946 673
rect 2893 602 2904 636
rect 2938 602 2946 636
rect 2893 565 2946 602
rect 2893 531 2904 565
rect 2938 531 2946 565
rect 2893 519 2946 531
<< mvndiffc >>
rect 42 156 76 190
rect 198 156 232 190
rect 1123 276 1157 310
rect 354 156 388 190
rect 497 132 531 166
rect 653 132 687 166
rect 813 132 847 166
rect 1111 121 1145 155
rect 1500 241 1534 275
rect 1500 149 1534 183
rect 1821 241 1855 275
rect 2284 228 2318 262
rect 2440 228 2474 262
rect 2565 228 2599 262
rect 2744 245 2778 279
rect 2744 145 2778 179
rect 2900 245 2934 279
rect 2900 145 2934 179
<< mvpdiffc >>
rect 39 697 73 731
rect 39 605 73 639
rect 195 701 229 735
rect 195 601 229 635
rect 351 697 385 731
rect 351 605 385 639
rect 1508 673 1542 707
rect 463 554 497 588
rect 673 554 707 588
rect 829 554 863 588
rect 1137 571 1171 605
rect 1329 554 1363 588
rect 1508 604 1542 638
rect 1508 535 1542 569
rect 1825 627 1859 661
rect 2276 684 2310 718
rect 2463 684 2497 718
rect 2748 673 2782 707
rect 2142 545 2176 579
rect 2298 527 2332 561
rect 2573 623 2607 657
rect 2573 531 2607 565
rect 2748 602 2782 636
rect 2748 531 2782 565
rect 2904 673 2938 707
rect 2904 602 2938 636
rect 2904 531 2938 565
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 2976 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
<< poly >>
rect 84 743 184 769
rect 240 743 340 769
rect 513 735 818 781
rect 1889 753 1989 773
rect 513 701 533 735
rect 567 701 818 735
rect 513 681 818 701
rect 562 613 662 639
rect 718 613 818 681
rect 876 707 982 735
rect 876 673 896 707
rect 930 673 982 707
rect 876 635 982 673
rect 882 613 982 635
rect 1024 695 1124 735
rect 1553 715 1653 741
rect 1695 715 1795 741
rect 1889 719 1915 753
rect 1949 719 1989 753
rect 2352 743 2452 769
rect 1024 661 1044 695
rect 1078 661 1124 695
rect 1024 613 1124 661
rect 1218 613 1318 639
rect 1374 613 1474 639
rect 84 533 184 593
rect 84 499 125 533
rect 159 499 184 533
rect 84 490 184 499
rect 84 465 187 490
rect 84 431 125 465
rect 159 431 187 465
rect 84 390 187 431
rect 240 390 340 593
rect 562 503 662 529
rect 497 413 662 503
rect 87 215 187 390
rect 232 370 343 390
rect 232 336 252 370
rect 286 336 343 370
rect 232 302 343 336
rect 232 268 252 302
rect 286 268 343 302
rect 232 241 343 268
rect 497 379 517 413
rect 551 403 662 413
rect 718 507 818 529
rect 718 447 840 507
rect 882 503 982 529
rect 718 417 946 447
rect 718 407 890 417
rect 551 379 597 403
rect 497 359 597 379
rect 840 383 890 407
rect 924 395 946 417
rect 1024 407 1124 529
rect 1218 503 1318 529
rect 924 383 958 395
rect 497 345 642 359
rect 497 311 517 345
rect 551 311 642 345
rect 497 259 642 311
rect 243 215 343 241
rect 542 191 642 259
rect 698 335 798 355
rect 698 301 743 335
rect 777 301 798 335
rect 698 267 798 301
rect 840 349 958 383
rect 840 315 890 349
rect 924 315 958 349
rect 1024 331 1100 407
rect 1168 357 1318 503
rect 1374 409 1474 529
rect 1889 599 1989 719
rect 2793 719 2893 745
rect 2618 669 2718 695
rect 2352 637 2452 659
rect 2031 599 2131 625
rect 2187 599 2287 625
rect 2352 592 2459 637
rect 2359 519 2459 592
rect 1553 493 1653 515
rect 1545 417 1653 493
rect 1695 493 1795 515
rect 1695 467 1847 493
rect 1889 489 1989 515
rect 1695 433 1742 467
rect 1776 447 1847 467
rect 1776 433 1989 447
rect 1695 417 1989 433
rect 1370 359 1503 409
rect 1168 335 1268 357
rect 840 295 958 315
rect 698 233 743 267
rect 777 233 798 267
rect 698 191 798 233
rect 858 191 958 295
rect 1000 311 1100 331
rect 1000 277 1043 311
rect 1077 277 1100 311
rect 1000 191 1100 277
rect 1370 325 1449 359
rect 1483 325 1503 359
rect 1370 309 1503 325
rect 1370 287 1470 309
rect 1545 287 1645 417
rect 1687 359 1757 375
rect 1687 325 1707 359
rect 1741 325 1757 359
rect 1799 355 1989 417
rect 1687 313 1757 325
rect 1687 287 1787 313
rect 1889 287 1989 355
rect 2031 427 2131 515
rect 2187 489 2287 515
rect 2359 497 2392 519
rect 2031 393 2077 427
rect 2111 393 2131 427
rect 2031 359 2131 393
rect 2031 325 2077 359
rect 2111 325 2131 359
rect 2031 287 2131 325
rect 2173 313 2287 489
rect 2329 485 2392 497
rect 2426 497 2459 519
rect 2618 497 2718 519
rect 2426 485 2718 497
rect 2793 493 2893 519
rect 2329 451 2718 485
rect 2329 417 2392 451
rect 2426 417 2718 451
rect 2329 397 2718 417
rect 2778 463 2893 493
rect 2778 429 2798 463
rect 2832 429 2893 463
rect 2173 287 2273 313
rect 2329 287 2429 397
rect 2610 287 2710 397
rect 2778 395 2893 429
rect 2778 361 2798 395
rect 2832 361 2893 395
rect 2778 313 2893 361
rect 2789 287 2889 313
rect 87 105 187 131
rect 243 105 343 131
rect 1168 171 1268 251
rect 1370 177 1470 203
rect 1168 137 1213 171
rect 1247 137 1268 171
rect 1889 177 1989 203
rect 2031 177 2131 203
rect 2173 161 2273 203
rect 2329 177 2429 203
rect 2610 177 2710 203
rect 1168 115 1268 137
rect 1545 115 1645 137
rect 542 81 642 107
rect 698 81 798 107
rect 858 81 958 107
rect 1000 81 1100 107
rect 1168 103 1645 115
rect 1687 111 1787 137
rect 2173 127 2193 161
rect 2227 127 2273 161
rect 1168 69 1213 103
rect 1247 69 1645 103
rect 2173 81 2273 127
rect 2789 111 2889 137
rect 1168 28 1645 69
<< polycont >>
rect 533 701 567 735
rect 896 673 930 707
rect 1915 719 1949 753
rect 1044 661 1078 695
rect 125 499 159 533
rect 125 431 159 465
rect 252 336 286 370
rect 252 268 286 302
rect 517 379 551 413
rect 890 383 924 417
rect 517 311 551 345
rect 743 301 777 335
rect 890 315 924 349
rect 1742 433 1776 467
rect 743 233 777 267
rect 1043 277 1077 311
rect 1449 325 1483 359
rect 1707 325 1741 359
rect 2077 393 2111 427
rect 2077 325 2111 359
rect 2392 485 2426 519
rect 2392 417 2426 451
rect 2798 429 2832 463
rect 2798 361 2832 395
rect 1213 137 1247 171
rect 2193 127 2227 161
rect 1213 69 1247 103
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 2976 831
rect 1739 753 1965 761
rect 23 731 73 747
rect 23 697 39 731
rect 23 639 73 697
rect 23 605 39 639
rect 23 293 73 605
rect 109 735 299 751
rect 109 701 115 735
rect 149 701 187 735
rect 229 701 259 735
rect 293 701 299 735
rect 109 635 299 701
rect 109 601 195 635
rect 229 601 299 635
rect 109 585 299 601
rect 335 731 401 747
rect 335 697 351 731
rect 385 697 401 731
rect 335 639 401 697
rect 335 605 351 639
rect 385 605 401 639
rect 335 589 401 605
rect 109 533 175 549
rect 109 499 125 533
rect 159 499 175 533
rect 109 465 175 499
rect 109 431 125 465
rect 159 431 175 465
rect 109 415 175 431
rect 338 489 401 589
rect 447 735 497 741
rect 447 701 453 735
rect 487 701 497 735
rect 447 588 497 701
rect 447 554 463 588
rect 447 525 497 554
rect 533 735 567 751
rect 1121 735 1187 741
rect 533 489 567 701
rect 338 455 567 489
rect 603 707 1001 723
rect 603 673 896 707
rect 930 673 1001 707
rect 603 657 1001 673
rect 236 370 302 379
rect 236 336 252 370
rect 286 336 302 370
rect 236 302 302 336
rect 236 293 252 302
rect 23 268 252 293
rect 286 268 302 302
rect 23 259 302 268
rect 23 190 76 259
rect 23 156 42 190
rect 23 123 76 156
rect 114 190 232 223
rect 114 156 198 190
rect 114 113 232 156
rect 114 79 120 113
rect 154 79 192 113
rect 226 79 232 113
rect 114 73 232 79
rect 268 87 302 259
rect 338 190 388 455
rect 501 413 567 419
rect 501 379 517 413
rect 551 379 567 413
rect 501 345 567 379
rect 501 311 517 345
rect 551 311 567 345
rect 501 305 567 311
rect 603 269 637 657
rect 338 156 354 190
rect 338 123 388 156
rect 424 235 637 269
rect 673 588 707 621
rect 424 87 458 235
rect 673 199 707 554
rect 743 335 777 657
rect 743 267 777 301
rect 743 217 777 233
rect 813 588 879 621
rect 813 554 829 588
rect 863 554 879 588
rect 813 521 879 554
rect 813 227 847 521
rect 967 465 1001 657
rect 1037 695 1085 711
rect 1037 661 1044 695
rect 1078 661 1085 695
rect 1037 535 1085 661
rect 1121 701 1127 735
rect 1161 701 1187 735
rect 1121 605 1187 701
rect 1415 735 1605 741
rect 1415 701 1421 735
rect 1455 701 1493 735
rect 1527 707 1565 735
rect 1542 701 1565 707
rect 1599 701 1605 735
rect 1415 673 1508 701
rect 1542 673 1605 701
rect 1415 638 1605 673
rect 1121 571 1137 605
rect 1171 571 1187 605
rect 1313 588 1379 621
rect 1313 569 1329 588
rect 1223 554 1329 569
rect 1363 554 1379 588
rect 1223 535 1379 554
rect 1415 604 1508 638
rect 1542 604 1605 638
rect 1415 569 1605 604
rect 1415 535 1508 569
rect 1542 535 1605 569
rect 1739 719 1915 753
rect 1949 719 1965 753
rect 2002 735 2192 741
rect 1739 569 1773 719
rect 2002 701 2008 735
rect 2042 701 2080 735
rect 2114 701 2152 735
rect 2186 701 2192 735
rect 1809 661 1932 683
rect 1809 627 1825 661
rect 1859 627 1932 661
rect 1809 605 1932 627
rect 1739 535 1862 569
rect 1037 501 1257 535
rect 1293 467 1792 499
rect 1293 465 1742 467
rect 883 417 931 433
rect 967 431 1327 465
rect 1726 433 1742 465
rect 1776 433 1792 467
rect 883 383 890 417
rect 924 395 931 417
rect 1363 395 1690 429
rect 1726 417 1792 433
rect 924 383 1397 395
rect 883 361 1397 383
rect 1656 375 1690 395
rect 1828 375 1862 535
rect 883 349 931 361
rect 1656 359 1862 375
rect 883 315 890 349
rect 924 315 931 349
rect 1433 325 1449 359
rect 1483 325 1620 359
rect 883 299 931 315
rect 1027 311 1173 325
rect 1433 311 1620 325
rect 1027 277 1043 311
rect 1077 310 1173 311
rect 1077 277 1123 310
rect 1027 276 1123 277
rect 1157 276 1173 310
rect 1027 263 1173 276
rect 1360 241 1500 275
rect 1534 241 1550 275
rect 268 53 458 87
rect 494 166 601 199
rect 494 132 497 166
rect 531 132 601 166
rect 494 113 601 132
rect 528 79 566 113
rect 600 79 601 113
rect 637 166 707 199
rect 637 132 653 166
rect 687 132 707 166
rect 637 99 707 132
rect 813 193 1263 227
rect 813 166 863 193
rect 847 132 863 166
rect 1197 171 1263 193
rect 813 99 863 132
rect 971 155 1161 157
rect 971 121 1111 155
rect 1145 121 1161 155
rect 971 113 1161 121
rect 494 73 601 79
rect 971 79 977 113
rect 1011 79 1049 113
rect 1083 79 1121 113
rect 1155 79 1161 113
rect 971 73 1161 79
rect 1197 137 1213 171
rect 1247 137 1263 171
rect 1197 103 1263 137
rect 1197 69 1213 103
rect 1247 69 1263 103
rect 1360 183 1550 241
rect 1360 149 1500 183
rect 1534 149 1550 183
rect 1586 202 1620 311
rect 1656 325 1707 359
rect 1741 341 1862 359
rect 1898 497 1932 605
rect 2002 579 2192 701
rect 2260 718 2310 751
rect 2260 684 2276 718
rect 2260 651 2310 684
rect 2346 735 2536 747
rect 2346 701 2352 735
rect 2386 701 2424 735
rect 2458 718 2496 735
rect 2458 701 2463 718
rect 2530 701 2536 735
rect 2346 684 2463 701
rect 2497 684 2536 701
rect 2346 671 2536 684
rect 2659 735 2848 741
rect 2659 701 2664 735
rect 2698 701 2736 735
rect 2770 707 2808 735
rect 2782 701 2808 707
rect 2842 701 2848 735
rect 2659 673 2748 701
rect 2782 673 2848 701
rect 2276 635 2310 651
rect 2573 657 2623 673
rect 2276 601 2512 635
rect 2002 545 2142 579
rect 2176 545 2192 579
rect 2002 533 2192 545
rect 2282 561 2348 565
rect 2282 527 2298 561
rect 2332 535 2348 561
rect 2332 527 2442 535
rect 2282 519 2442 527
rect 2282 497 2392 519
rect 1898 485 2392 497
rect 2426 485 2442 519
rect 1898 463 2442 485
rect 1741 325 1757 341
rect 1656 309 1757 325
rect 1898 295 1932 463
rect 2376 451 2442 463
rect 2061 393 2077 427
rect 2111 393 2127 427
rect 2376 417 2392 451
rect 2426 417 2442 451
rect 2376 401 2442 417
rect 2061 365 2127 393
rect 2478 365 2512 601
rect 2061 359 2512 365
rect 2061 325 2077 359
rect 2111 331 2512 359
rect 2607 623 2623 657
rect 2573 565 2623 623
rect 2607 531 2623 565
rect 2573 479 2623 531
rect 2659 636 2848 673
rect 2659 602 2748 636
rect 2782 602 2848 636
rect 2659 565 2848 602
rect 2659 531 2748 565
rect 2782 531 2848 565
rect 2659 515 2848 531
rect 2884 707 2954 723
rect 2884 673 2904 707
rect 2938 673 2954 707
rect 2884 636 2954 673
rect 2884 602 2904 636
rect 2938 602 2954 636
rect 2884 565 2954 602
rect 2884 531 2904 565
rect 2938 531 2954 565
rect 2573 463 2848 479
rect 2573 445 2798 463
rect 2111 325 2127 331
rect 2061 309 2127 325
rect 1805 275 1932 295
rect 1805 241 1821 275
rect 1855 241 1932 275
rect 1805 238 1932 241
rect 2268 262 2386 295
rect 2268 228 2284 262
rect 2318 228 2386 262
rect 2177 202 2232 208
rect 1586 168 2232 202
rect 1360 113 1550 149
rect 1360 79 1366 113
rect 1400 79 1438 113
rect 1472 79 1510 113
rect 1544 79 1550 113
rect 1657 161 2232 168
rect 1657 127 2193 161
rect 2227 127 2232 161
rect 1657 111 2232 127
rect 2268 113 2386 228
rect 2424 262 2490 331
rect 2573 295 2615 445
rect 2782 429 2798 445
rect 2832 429 2848 463
rect 2782 395 2848 429
rect 2782 361 2798 395
rect 2832 361 2848 395
rect 2782 345 2848 361
rect 2424 228 2440 262
rect 2474 228 2490 262
rect 2424 195 2490 228
rect 2549 262 2615 295
rect 2549 228 2565 262
rect 2599 228 2615 262
rect 2549 195 2615 228
rect 2651 279 2841 295
rect 2651 245 2744 279
rect 2778 245 2841 279
rect 1360 73 1550 79
rect 2268 79 2274 113
rect 2308 79 2346 113
rect 2380 79 2386 113
rect 2268 73 2386 79
rect 2651 179 2841 245
rect 2651 145 2744 179
rect 2778 145 2841 179
rect 2651 113 2841 145
rect 2884 279 2954 531
rect 2884 245 2900 279
rect 2934 245 2954 279
rect 2884 179 2954 245
rect 2884 145 2900 179
rect 2934 145 2954 179
rect 2884 129 2954 145
rect 2651 79 2657 113
rect 2691 79 2729 113
rect 2763 79 2801 113
rect 2835 79 2841 113
rect 2651 73 2841 79
rect 1197 53 1263 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 115 701 149 735
rect 187 701 195 735
rect 195 701 221 735
rect 259 701 293 735
rect 453 701 487 735
rect 120 79 154 113
rect 192 79 226 113
rect 1127 701 1161 735
rect 1421 701 1455 735
rect 1493 707 1527 735
rect 1493 701 1508 707
rect 1508 701 1527 707
rect 1565 701 1599 735
rect 2008 701 2042 735
rect 2080 701 2114 735
rect 2152 701 2186 735
rect 494 79 528 113
rect 566 79 600 113
rect 977 79 1011 113
rect 1049 79 1083 113
rect 1121 79 1155 113
rect 2352 701 2386 735
rect 2424 701 2458 735
rect 2496 718 2530 735
rect 2496 701 2497 718
rect 2497 701 2530 718
rect 2664 701 2698 735
rect 2736 707 2770 735
rect 2736 701 2748 707
rect 2748 701 2770 707
rect 2808 701 2842 735
rect 1366 79 1400 113
rect 1438 79 1472 113
rect 1510 79 1544 113
rect 2274 79 2308 113
rect 2346 79 2380 113
rect 2657 79 2691 113
rect 2729 79 2763 113
rect 2801 79 2835 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< metal1 >>
rect 0 831 2976 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 2976 831
rect 0 791 2976 797
rect 0 735 2976 763
rect 0 701 115 735
rect 149 701 187 735
rect 221 701 259 735
rect 293 701 453 735
rect 487 701 1127 735
rect 1161 701 1421 735
rect 1455 701 1493 735
rect 1527 701 1565 735
rect 1599 701 2008 735
rect 2042 701 2080 735
rect 2114 701 2152 735
rect 2186 701 2352 735
rect 2386 701 2424 735
rect 2458 701 2496 735
rect 2530 701 2664 735
rect 2698 701 2736 735
rect 2770 701 2808 735
rect 2842 701 2976 735
rect 0 689 2976 701
rect 0 113 2976 125
rect 0 79 120 113
rect 154 79 192 113
rect 226 79 494 113
rect 528 79 566 113
rect 600 79 977 113
rect 1011 79 1049 113
rect 1083 79 1121 113
rect 1155 79 1366 113
rect 1400 79 1438 113
rect 1472 79 1510 113
rect 1544 79 2274 113
rect 2308 79 2346 113
rect 2380 79 2657 113
rect 2691 79 2729 113
rect 2763 79 2801 113
rect 2835 79 2976 113
rect 0 51 2976 79
rect 0 17 2976 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
rect 0 -23 2976 -17
<< labels >>
flabel comment s 1059 477 1059 477 0 FreeSans 200 90 0 0 no_jumper_check
flabel comment s 687 739 687 739 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfstp_1
flabel metal1 s 0 51 2976 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 0 2976 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 689 2976 763 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 791 2976 814 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 1663 168 1697 202 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1759 168 1793 202 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1855 168 1889 202 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1951 168 1985 202 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 2047 168 2081 202 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 2143 168 2177 202 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2911 168 2945 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2911 242 2945 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2911 316 2945 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2911 390 2945 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2911 464 2945 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2911 538 2945 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2911 612 2945 646 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
rlabel locali s 2268 73 2386 295 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 2651 73 2841 295 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 494 73 601 199 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 971 73 1161 157 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 1360 73 1550 275 1 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 51 2976 125 1 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 -23 2976 23 1 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 791 2976 837 1 VPB
port 6 nsew power bidirectional
rlabel locali s 2002 533 2192 741 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2346 671 2536 747 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2659 515 2848 741 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 447 525 497 741 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 1121 571 1187 741 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 1415 535 1605 741 1 VPWR
port 7 nsew power bidirectional
rlabel metal1 s 0 689 2976 763 1 VPWR
port 7 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 2976 814
string GDS_END 918942
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 889776
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
