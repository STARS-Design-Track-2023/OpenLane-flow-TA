magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__hvdfl1sd2__example_55959141808316  sky130_fd_pr__hvdfl1sd2__example_55959141808316_0
timestamp 1686671242
transform 1 0 132 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808137  sky130_fd_pr__hvdfl1sd__example_55959141808137_0
timestamp 1686671242
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808506  sky130_fd_pr__hvdftpl1s2__example_55959141808506_0
timestamp 1686671242
transform 1 0 320 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 48481298
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48479596
<< end >>
