magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect 2713 184 3247 456
<< pwell >>
rect 54 955 306 2661
rect 72 861 306 955
rect 72 10 424 861
rect 610 10 962 424
<< mvnmos >>
rect 98 682 398 782
rect 98 526 398 626
rect 98 245 398 345
rect 98 89 398 189
rect 636 245 936 345
rect 636 89 936 189
<< mvpmos >>
rect 2832 250 2952 390
rect 3008 250 3128 390
<< mvnnmos >>
rect 80 1863 280 2043
rect 80 1627 280 1807
rect 80 1270 280 1450
rect 80 1034 280 1214
<< nmoslvt >>
rect 80 2552 280 2582
rect 80 2466 280 2496
rect 80 2380 280 2410
rect 80 2294 280 2324
<< ndiff >>
rect 80 2627 280 2635
rect 80 2593 92 2627
rect 126 2593 160 2627
rect 194 2593 228 2627
rect 262 2593 280 2627
rect 80 2582 280 2593
rect 80 2541 280 2552
rect 80 2507 92 2541
rect 126 2507 160 2541
rect 194 2507 228 2541
rect 262 2507 280 2541
rect 80 2496 280 2507
rect 80 2455 280 2466
rect 80 2421 92 2455
rect 126 2421 160 2455
rect 194 2421 228 2455
rect 262 2421 280 2455
rect 80 2410 280 2421
rect 80 2369 280 2380
rect 80 2335 92 2369
rect 126 2335 160 2369
rect 194 2335 228 2369
rect 262 2335 280 2369
rect 80 2324 280 2335
rect 80 2283 280 2294
rect 80 2249 92 2283
rect 126 2249 160 2283
rect 194 2249 228 2283
rect 262 2249 280 2283
rect 80 2241 280 2249
<< mvndiff >>
rect 80 2088 280 2096
rect 80 2054 92 2088
rect 126 2054 160 2088
rect 194 2054 228 2088
rect 262 2054 280 2088
rect 80 2043 280 2054
rect 80 1852 280 1863
rect 80 1818 92 1852
rect 126 1818 160 1852
rect 194 1818 228 1852
rect 262 1818 280 1852
rect 80 1807 280 1818
rect 80 1616 280 1627
rect 80 1582 92 1616
rect 126 1582 160 1616
rect 194 1582 228 1616
rect 262 1582 280 1616
rect 80 1574 280 1582
rect 80 1495 280 1503
rect 80 1461 98 1495
rect 132 1461 166 1495
rect 200 1461 234 1495
rect 268 1461 280 1495
rect 80 1450 280 1461
rect 80 1259 280 1270
rect 80 1225 98 1259
rect 132 1225 166 1259
rect 200 1225 234 1259
rect 268 1225 280 1259
rect 80 1214 280 1225
rect 80 1023 280 1034
rect 80 989 98 1023
rect 132 989 166 1023
rect 200 989 234 1023
rect 268 989 280 1023
rect 80 981 280 989
rect 98 827 398 835
rect 98 793 110 827
rect 144 793 178 827
rect 212 793 246 827
rect 280 793 314 827
rect 348 793 398 827
rect 98 782 398 793
rect 98 671 398 682
rect 98 637 110 671
rect 144 637 178 671
rect 212 637 246 671
rect 280 637 314 671
rect 348 637 398 671
rect 98 626 398 637
rect 98 515 398 526
rect 98 481 110 515
rect 144 481 178 515
rect 212 481 246 515
rect 280 481 314 515
rect 348 481 398 515
rect 98 473 398 481
rect 98 390 398 398
rect 98 356 110 390
rect 144 356 178 390
rect 212 356 246 390
rect 280 356 314 390
rect 348 356 398 390
rect 98 345 398 356
rect 636 390 936 398
rect 636 356 648 390
rect 682 356 716 390
rect 750 356 784 390
rect 818 356 852 390
rect 886 356 936 390
rect 636 345 936 356
rect 98 234 398 245
rect 98 200 110 234
rect 144 200 178 234
rect 212 200 246 234
rect 280 200 314 234
rect 348 200 398 234
rect 98 189 398 200
rect 636 234 936 245
rect 636 200 648 234
rect 682 200 716 234
rect 750 200 784 234
rect 818 200 852 234
rect 886 200 936 234
rect 636 189 936 200
rect 98 78 398 89
rect 98 44 110 78
rect 144 44 178 78
rect 212 44 246 78
rect 280 44 314 78
rect 348 44 398 78
rect 98 36 398 44
rect 636 78 936 89
rect 636 44 648 78
rect 682 44 716 78
rect 750 44 784 78
rect 818 44 852 78
rect 886 44 936 78
rect 636 36 936 44
<< mvpdiff >>
rect 2779 364 2832 390
rect 2779 330 2787 364
rect 2821 330 2832 364
rect 2779 296 2832 330
rect 2779 262 2787 296
rect 2821 262 2832 296
rect 2779 250 2832 262
rect 2952 364 3008 390
rect 2952 330 2963 364
rect 2997 330 3008 364
rect 2952 296 3008 330
rect 2952 262 2963 296
rect 2997 262 3008 296
rect 2952 250 3008 262
rect 3128 364 3181 390
rect 3128 330 3139 364
rect 3173 330 3181 364
rect 3128 296 3181 330
rect 3128 262 3139 296
rect 3173 262 3181 296
rect 3128 250 3181 262
<< ndiffc >>
rect 92 2593 126 2627
rect 160 2593 194 2627
rect 228 2593 262 2627
rect 92 2507 126 2541
rect 160 2507 194 2541
rect 228 2507 262 2541
rect 92 2421 126 2455
rect 160 2421 194 2455
rect 228 2421 262 2455
rect 92 2335 126 2369
rect 160 2335 194 2369
rect 228 2335 262 2369
rect 92 2249 126 2283
rect 160 2249 194 2283
rect 228 2249 262 2283
<< mvndiffc >>
rect 92 2054 126 2088
rect 160 2054 194 2088
rect 228 2054 262 2088
rect 92 1818 126 1852
rect 160 1818 194 1852
rect 228 1818 262 1852
rect 92 1582 126 1616
rect 160 1582 194 1616
rect 228 1582 262 1616
rect 98 1461 132 1495
rect 166 1461 200 1495
rect 234 1461 268 1495
rect 98 1225 132 1259
rect 166 1225 200 1259
rect 234 1225 268 1259
rect 98 989 132 1023
rect 166 989 200 1023
rect 234 989 268 1023
rect 110 793 144 827
rect 178 793 212 827
rect 246 793 280 827
rect 314 793 348 827
rect 110 637 144 671
rect 178 637 212 671
rect 246 637 280 671
rect 314 637 348 671
rect 110 481 144 515
rect 178 481 212 515
rect 246 481 280 515
rect 314 481 348 515
rect 110 356 144 390
rect 178 356 212 390
rect 246 356 280 390
rect 314 356 348 390
rect 648 356 682 390
rect 716 356 750 390
rect 784 356 818 390
rect 852 356 886 390
rect 110 200 144 234
rect 178 200 212 234
rect 246 200 280 234
rect 314 200 348 234
rect 648 200 682 234
rect 716 200 750 234
rect 784 200 818 234
rect 852 200 886 234
rect 110 44 144 78
rect 178 44 212 78
rect 246 44 280 78
rect 314 44 348 78
rect 648 44 682 78
rect 716 44 750 78
rect 784 44 818 78
rect 852 44 886 78
<< mvpdiffc >>
rect 2787 330 2821 364
rect 2787 262 2821 296
rect 2963 330 2997 364
rect 2963 262 2997 296
rect 3139 330 3173 364
rect 3139 262 3173 296
<< poly >>
rect 312 2584 378 2600
rect 312 2582 328 2584
rect 48 2552 80 2582
rect 280 2552 328 2582
rect 312 2550 328 2552
rect 362 2550 378 2584
rect 312 2516 378 2550
rect 312 2496 328 2516
rect 48 2466 80 2496
rect 280 2482 328 2496
rect 362 2482 378 2516
rect 280 2466 378 2482
rect 48 2380 80 2410
rect 280 2394 378 2410
rect 280 2380 328 2394
rect 312 2360 328 2380
rect 362 2360 378 2394
rect 312 2326 378 2360
rect 312 2324 328 2326
rect 48 2294 80 2324
rect 280 2294 328 2324
rect 312 2292 328 2294
rect 362 2292 378 2326
rect 312 2276 378 2292
rect 48 1863 80 2043
rect 280 2027 378 2043
rect 280 1993 328 2027
rect 362 1993 378 2027
rect 280 1954 378 1993
rect 280 1920 328 1954
rect 362 1920 378 1954
rect 280 1881 378 1920
rect 280 1863 328 1881
rect 312 1847 328 1863
rect 362 1847 378 1881
rect 312 1808 378 1847
rect 312 1807 328 1808
rect 48 1627 80 1807
rect 280 1774 328 1807
rect 362 1774 378 1808
rect 280 1735 378 1774
rect 280 1701 328 1735
rect 362 1701 378 1735
rect 280 1662 378 1701
rect 280 1628 328 1662
rect 362 1628 378 1662
rect 280 1627 378 1628
rect 312 1589 378 1627
rect 312 1555 328 1589
rect 362 1555 378 1589
rect 312 1516 378 1555
rect 312 1482 328 1516
rect 362 1482 378 1516
rect 312 1450 378 1482
rect 48 1270 80 1450
rect 280 1444 378 1450
rect 280 1410 328 1444
rect 362 1410 378 1444
rect 280 1372 378 1410
rect 280 1338 328 1372
rect 362 1338 378 1372
rect 280 1300 378 1338
rect 280 1270 328 1300
rect 312 1266 328 1270
rect 362 1266 378 1300
rect 312 1228 378 1266
rect 312 1214 328 1228
rect 48 1034 80 1214
rect 280 1194 328 1214
rect 362 1194 378 1228
rect 280 1156 378 1194
rect 280 1122 328 1156
rect 362 1122 378 1156
rect 280 1084 378 1122
rect 280 1050 328 1084
rect 362 1050 378 1084
rect 280 1034 378 1050
rect 66 682 98 782
rect 398 766 496 782
rect 398 732 446 766
rect 480 732 496 766
rect 398 682 496 732
rect 430 671 496 682
rect 430 637 446 671
rect 480 637 496 671
rect 430 626 496 637
rect 66 526 98 626
rect 398 576 496 626
rect 398 542 446 576
rect 480 542 496 576
rect 398 526 496 542
rect 2813 472 2952 488
rect 2813 438 2829 472
rect 2863 438 2902 472
rect 2936 438 2952 472
rect 2813 422 2952 438
rect 2832 390 2952 422
rect 3008 472 3147 488
rect 3008 438 3024 472
rect 3058 438 3097 472
rect 3131 438 3147 472
rect 3008 422 3147 438
rect 3008 390 3128 422
rect 66 245 98 345
rect 398 329 496 345
rect 398 295 446 329
rect 480 295 496 329
rect 398 245 496 295
rect 430 234 496 245
rect 430 200 446 234
rect 480 200 496 234
rect 430 189 496 200
rect 66 89 98 189
rect 398 139 496 189
rect 398 105 446 139
rect 480 105 496 139
rect 398 89 496 105
rect 538 329 636 345
rect 538 295 554 329
rect 588 295 636 329
rect 538 245 636 295
rect 936 245 968 345
rect 538 234 604 245
rect 538 200 554 234
rect 588 200 604 234
rect 538 189 604 200
rect 2832 218 2952 250
rect 3008 218 3128 250
rect 538 139 636 189
rect 538 105 554 139
rect 588 105 636 139
rect 538 89 636 105
rect 936 89 968 189
<< polycont >>
rect 328 2550 362 2584
rect 328 2482 362 2516
rect 328 2360 362 2394
rect 328 2292 362 2326
rect 328 1993 362 2027
rect 328 1920 362 1954
rect 328 1847 362 1881
rect 328 1774 362 1808
rect 328 1701 362 1735
rect 328 1628 362 1662
rect 328 1555 362 1589
rect 328 1482 362 1516
rect 328 1410 362 1444
rect 328 1338 362 1372
rect 328 1266 362 1300
rect 328 1194 362 1228
rect 328 1122 362 1156
rect 328 1050 362 1084
rect 446 732 480 766
rect 446 637 480 671
rect 446 542 480 576
rect 2829 438 2863 472
rect 2902 438 2936 472
rect 3024 438 3058 472
rect 3097 438 3131 472
rect 446 295 480 329
rect 446 200 480 234
rect 446 105 480 139
rect 554 295 588 329
rect 554 200 588 234
rect 554 105 588 139
<< locali >>
rect -31 2627 278 2649
rect -31 2593 92 2627
rect 126 2593 160 2627
rect 194 2593 228 2627
rect 262 2593 278 2627
rect 328 2588 362 2600
rect 76 2539 92 2541
rect 76 2507 88 2539
rect 126 2507 160 2541
rect 194 2507 228 2541
rect 262 2507 278 2541
rect 328 2516 362 2550
rect 122 2505 160 2507
rect 328 2466 362 2478
rect -31 2455 278 2466
rect -31 2421 92 2455
rect 126 2421 160 2455
rect 194 2421 228 2455
rect 262 2421 278 2455
rect -31 2410 278 2421
rect 328 2398 362 2410
rect 328 2394 334 2398
rect 214 2369 252 2370
rect 76 2335 92 2369
rect 126 2335 160 2369
rect 214 2336 228 2369
rect 362 2360 368 2364
rect 194 2335 228 2336
rect 262 2335 278 2336
rect 328 2326 368 2360
rect 362 2322 368 2326
rect -31 2283 278 2291
rect -31 2249 92 2283
rect 126 2249 160 2283
rect 194 2249 228 2283
rect 262 2249 278 2283
rect 328 2288 334 2292
rect 328 2276 362 2288
rect -31 2235 278 2249
rect 76 2054 92 2088
rect 126 2054 160 2088
rect 200 2084 228 2088
rect 194 2054 228 2084
rect 262 2054 278 2088
rect 166 2046 200 2054
rect 328 2031 362 2043
rect 328 2027 334 2031
rect 362 1993 368 1997
rect 328 1958 368 1993
rect 328 1954 334 1958
rect 362 1920 368 1924
rect 328 1885 368 1920
rect 76 1818 92 1852
rect 126 1818 160 1852
rect 194 1818 228 1852
rect 262 1818 292 1850
rect 258 1812 292 1818
rect 328 1881 334 1885
rect 362 1847 368 1851
rect 328 1812 368 1847
rect 328 1808 334 1812
rect 362 1774 368 1778
rect 328 1739 368 1774
rect 328 1735 334 1739
rect 362 1701 368 1705
rect 166 1616 200 1634
rect 328 1666 368 1701
rect 328 1662 334 1666
rect 362 1628 368 1632
rect 76 1582 92 1616
rect 126 1582 160 1616
rect 194 1596 228 1616
rect 200 1582 228 1596
rect 262 1582 278 1616
rect 328 1593 368 1628
rect 328 1589 334 1593
rect 362 1555 368 1559
rect 328 1520 368 1555
rect 82 1461 98 1495
rect 132 1461 166 1495
rect 200 1461 234 1495
rect 268 1461 292 1484
rect 258 1446 292 1461
rect 328 1516 334 1520
rect 362 1482 368 1486
rect 328 1447 368 1482
rect 328 1444 334 1447
rect 362 1410 368 1413
rect 328 1374 368 1410
rect 328 1372 334 1374
rect 362 1338 368 1340
rect 328 1301 368 1338
rect 328 1300 334 1301
rect 362 1266 368 1267
rect 82 1258 84 1259
rect 82 1225 98 1258
rect 132 1225 166 1259
rect 200 1225 234 1259
rect 268 1225 284 1259
rect 328 1228 368 1266
rect 362 1227 368 1228
rect 84 1220 118 1225
rect 328 1193 334 1194
rect 328 1156 368 1193
rect 362 1153 368 1156
rect 328 1119 334 1122
rect 258 1023 292 1061
rect 328 1084 368 1119
rect 362 1079 368 1084
rect 328 1045 334 1050
rect 328 1034 362 1045
rect 82 989 98 1023
rect 132 989 166 1023
rect 200 989 234 1023
rect 94 793 110 827
rect 144 793 178 827
rect 212 793 246 827
rect 280 793 314 827
rect 348 793 370 794
rect 336 756 370 793
rect 446 770 480 782
rect 446 671 480 732
rect 94 637 110 671
rect 144 637 178 671
rect 212 637 246 671
rect 280 637 314 671
rect 348 637 364 671
rect 166 633 200 637
rect 446 576 480 637
rect 446 526 480 538
rect 94 481 110 515
rect 144 481 178 515
rect 212 481 246 515
rect 280 481 314 515
rect 348 481 370 515
rect 336 477 370 481
rect 2859 472 2906 473
rect 3021 472 3055 490
rect 2813 439 2825 472
rect 2813 438 2829 439
rect 2863 438 2902 472
rect 2940 439 2952 472
rect 2936 438 2952 439
rect 3008 443 3024 472
rect 3008 438 3021 443
rect 3058 438 3097 472
rect 3131 438 3147 472
rect 167 390 201 392
rect 94 356 110 390
rect 144 356 178 390
rect 212 356 246 390
rect 280 356 314 390
rect 348 356 364 390
rect 632 356 648 390
rect 682 356 716 390
rect 750 356 784 390
rect 818 356 852 390
rect 886 356 902 390
rect 2787 369 2821 380
rect 167 354 201 356
rect 446 333 480 345
rect 446 234 480 295
rect 94 200 110 234
rect 144 200 178 234
rect 212 200 246 234
rect 280 200 314 234
rect 348 200 364 234
rect 258 196 292 200
rect 446 139 480 200
rect 446 89 480 101
rect 554 333 588 345
rect 554 234 588 295
rect 2787 297 2821 330
rect 2787 246 2821 262
rect 2963 364 2997 380
rect 2963 296 2997 330
rect 2963 246 2997 262
rect 3139 369 3173 380
rect 3139 364 3159 369
rect 3173 330 3193 335
rect 3139 297 3193 330
rect 3139 296 3159 297
rect 3139 246 3173 262
rect 632 200 644 234
rect 682 200 716 234
rect 750 200 780 234
rect 818 200 852 234
rect 886 200 902 234
rect 554 139 588 200
rect 554 89 588 101
rect 167 78 201 80
rect 94 44 110 78
rect 144 44 178 78
rect 212 44 246 78
rect 280 44 314 78
rect 348 44 364 78
rect 632 44 648 78
rect 682 44 716 78
rect 750 44 784 78
rect 818 44 852 78
rect 886 44 902 78
rect 167 42 201 44
<< viali >>
rect 328 2584 362 2588
rect 328 2554 362 2584
rect 88 2507 92 2539
rect 92 2507 122 2539
rect 160 2507 194 2539
rect 88 2505 122 2507
rect 160 2505 194 2507
rect 328 2482 362 2512
rect 328 2478 362 2482
rect 334 2394 368 2398
rect 180 2369 214 2370
rect 252 2369 286 2370
rect 180 2336 194 2369
rect 194 2336 214 2369
rect 252 2336 262 2369
rect 262 2336 286 2369
rect 334 2364 362 2394
rect 362 2364 368 2394
rect 334 2292 362 2322
rect 362 2292 368 2322
rect 334 2288 368 2292
rect 166 2088 200 2118
rect 166 2084 194 2088
rect 194 2084 200 2088
rect 166 2012 200 2046
rect 334 2027 368 2031
rect 334 1997 362 2027
rect 362 1997 368 2027
rect 334 1954 368 1958
rect 334 1924 362 1954
rect 362 1924 368 1954
rect 258 1852 292 1884
rect 258 1850 262 1852
rect 262 1850 292 1852
rect 258 1778 292 1812
rect 334 1881 368 1885
rect 334 1851 362 1881
rect 362 1851 368 1881
rect 334 1808 368 1812
rect 334 1778 362 1808
rect 362 1778 368 1808
rect 334 1735 368 1739
rect 334 1705 362 1735
rect 362 1705 368 1735
rect 166 1634 200 1668
rect 334 1662 368 1666
rect 334 1632 362 1662
rect 362 1632 368 1662
rect 166 1582 194 1596
rect 194 1582 200 1596
rect 334 1589 368 1593
rect 166 1562 200 1582
rect 334 1559 362 1589
rect 362 1559 368 1589
rect 258 1495 292 1518
rect 258 1484 268 1495
rect 268 1484 292 1495
rect 258 1412 292 1446
rect 334 1516 368 1520
rect 334 1486 362 1516
rect 362 1486 368 1516
rect 334 1444 368 1447
rect 334 1413 362 1444
rect 362 1413 368 1444
rect 334 1372 368 1374
rect 334 1340 362 1372
rect 362 1340 368 1372
rect 334 1300 368 1301
rect 84 1259 118 1292
rect 334 1267 362 1300
rect 362 1267 368 1300
rect 84 1258 98 1259
rect 98 1258 118 1259
rect 84 1186 118 1220
rect 334 1194 362 1227
rect 362 1194 368 1227
rect 334 1193 368 1194
rect 334 1122 362 1153
rect 362 1122 368 1153
rect 334 1119 368 1122
rect 258 1061 292 1095
rect 334 1050 362 1079
rect 362 1050 368 1079
rect 334 1045 368 1050
rect 258 989 268 1023
rect 268 989 292 1023
rect 336 827 370 828
rect 336 794 348 827
rect 348 794 370 827
rect 336 722 370 756
rect 446 766 480 770
rect 446 736 480 766
rect 166 671 200 705
rect 446 637 480 671
rect 166 599 200 633
rect 336 515 370 549
rect 446 542 480 572
rect 446 538 480 542
rect 336 443 370 477
rect 3021 490 3055 524
rect 2825 472 2859 473
rect 2906 472 2940 473
rect 2825 439 2829 472
rect 2829 439 2859 472
rect 2906 439 2936 472
rect 2936 439 2940 472
rect 3021 438 3024 443
rect 3024 438 3055 443
rect 167 392 201 426
rect 3021 409 3055 438
rect 2787 364 2821 369
rect 167 320 201 354
rect 446 329 480 333
rect 446 299 480 329
rect 258 234 292 268
rect 446 200 480 234
rect 258 162 292 196
rect 167 80 201 114
rect 446 105 480 135
rect 446 101 480 105
rect 554 329 588 333
rect 554 299 588 329
rect 2787 335 2821 364
rect 2787 296 2821 297
rect 2787 263 2821 296
rect 3159 364 3193 369
rect 3159 335 3173 364
rect 3173 335 3193 364
rect 3159 296 3193 297
rect 3159 263 3173 296
rect 3173 263 3193 296
rect 554 200 588 234
rect 644 200 648 234
rect 648 200 678 234
rect 780 200 784 234
rect 784 200 814 234
rect 554 105 588 135
rect 554 101 588 105
rect 167 8 201 42
<< metal1 >>
rect 322 2588 368 2600
rect 322 2554 328 2588
rect 362 2554 368 2588
rect 76 2539 206 2545
rect 76 2505 88 2539
rect 122 2505 160 2539
rect 194 2505 206 2539
rect 76 2499 206 2505
rect 322 2512 368 2554
rect 78 1292 124 2499
rect 322 2478 328 2512
rect 362 2478 368 2512
rect 322 2466 368 2478
rect 328 2398 374 2410
rect 168 2370 298 2376
rect 168 2336 180 2370
rect 214 2336 252 2370
rect 286 2336 298 2370
rect 168 2330 298 2336
rect 78 1258 84 1292
rect 118 1258 124 1292
rect 78 1220 124 1258
rect 78 1186 84 1220
rect 118 1186 124 1220
rect 78 1174 124 1186
rect 160 2118 206 2130
rect 160 2084 166 2118
rect 200 2084 206 2118
rect 160 2046 206 2084
rect 160 2012 166 2046
rect 200 2012 206 2046
rect 160 1668 206 2012
rect 252 1884 298 2330
rect 328 2364 334 2398
rect 368 2364 374 2398
rect 328 2322 374 2364
rect 328 2288 334 2322
rect 368 2288 374 2322
rect 328 2276 374 2288
rect 252 1850 258 1884
rect 292 1850 298 1884
rect 252 1812 298 1850
rect 252 1778 258 1812
rect 292 1778 298 1812
rect 252 1766 298 1778
rect 328 2031 374 2043
rect 328 1997 334 2031
rect 368 1997 374 2031
rect 328 1958 374 1997
rect 328 1924 334 1958
rect 368 1924 374 1958
rect 328 1885 374 1924
rect 328 1851 334 1885
rect 368 1851 374 1885
rect 328 1812 374 1851
rect 328 1778 334 1812
rect 368 1778 374 1812
rect 160 1634 166 1668
rect 200 1634 206 1668
rect 160 1596 206 1634
rect 160 1562 166 1596
rect 200 1562 206 1596
rect 160 705 206 1562
rect 328 1739 374 1778
rect 328 1705 334 1739
rect 368 1705 374 1739
rect 328 1666 374 1705
rect 328 1632 334 1666
rect 368 1632 374 1666
rect 328 1593 374 1632
rect 328 1559 334 1593
rect 368 1559 374 1593
rect 160 671 166 705
rect 200 671 206 705
rect 160 633 206 671
rect 160 599 166 633
rect 200 599 206 633
rect 160 587 206 599
rect 252 1518 298 1530
rect 252 1484 258 1518
rect 292 1484 298 1518
rect 252 1446 298 1484
rect 252 1412 258 1446
rect 292 1412 298 1446
rect 252 1095 298 1412
rect 252 1061 258 1095
rect 292 1061 298 1095
rect 252 1023 298 1061
rect 328 1520 374 1559
rect 328 1486 334 1520
rect 368 1486 374 1520
rect 328 1447 374 1486
rect 328 1413 334 1447
rect 368 1413 374 1447
rect 328 1374 374 1413
rect 328 1340 334 1374
rect 368 1340 374 1374
rect 328 1301 374 1340
rect 328 1267 334 1301
rect 368 1267 374 1301
rect 328 1227 374 1267
rect 328 1193 334 1227
rect 368 1193 374 1227
rect 328 1153 374 1193
rect 328 1119 334 1153
rect 368 1119 374 1153
rect 328 1079 374 1119
rect 328 1045 334 1079
rect 368 1045 374 1079
rect 328 1033 374 1045
rect 252 989 258 1023
rect 292 989 298 1023
rect 161 426 207 438
rect 161 392 167 426
rect 201 392 207 426
rect 161 354 207 392
rect 161 349 167 354
rect 79 297 85 349
rect 137 297 149 349
rect 201 297 207 354
rect 161 114 207 297
rect 252 268 298 989
rect 330 794 336 872
rect 388 820 400 872
rect 452 820 458 872
rect 3047 820 3053 872
rect 3105 820 3117 872
rect 3169 820 3199 872
rect 370 794 376 820
rect 330 756 376 794
rect 330 722 336 756
rect 370 722 376 756
rect 330 549 376 722
rect 330 515 336 549
rect 370 515 376 549
rect 330 477 376 515
rect 330 443 336 477
rect 370 443 376 477
rect 330 430 376 443
rect 440 770 486 782
rect 440 736 446 770
rect 480 736 486 770
rect 440 671 486 736
rect 440 637 446 671
rect 480 637 486 671
rect 440 572 486 637
rect 440 538 446 572
rect 480 538 486 572
rect 252 234 258 268
rect 292 234 298 268
rect 252 196 298 234
rect 252 162 258 196
rect 292 162 298 196
rect 252 150 298 162
rect 440 333 486 538
rect 3015 524 3061 536
rect 3015 490 3021 524
rect 3055 490 3061 524
rect 2813 473 2952 479
rect 2813 439 2825 473
rect 2859 439 2906 473
rect 2940 439 2952 473
rect 2813 433 2952 439
rect 3015 443 3061 490
rect 3015 425 3021 443
rect 3009 419 3021 425
rect 3055 419 3061 443
rect 2781 369 2827 381
tri 2827 369 2839 381 sw
rect 440 299 446 333
rect 480 299 486 333
rect 440 234 486 299
rect 440 200 446 234
rect 480 200 486 234
rect 161 80 167 114
rect 201 80 207 114
rect 440 135 486 200
rect 440 101 446 135
rect 480 101 486 135
rect 440 89 486 101
rect 548 333 594 345
rect 548 299 554 333
rect 588 299 594 333
rect 548 234 594 299
rect 548 200 554 234
rect 588 200 594 234
rect 548 135 594 200
rect 632 297 638 349
rect 690 297 703 349
rect 755 297 768 349
rect 820 297 826 349
rect 632 234 826 297
rect 2781 263 2787 369
rect 2821 349 2839 369
tri 2839 349 2859 369 sw
rect 3009 355 3061 367
rect 2839 297 2851 349
rect 2903 297 2909 349
rect 3009 297 3061 303
rect 3153 369 3199 820
rect 3153 335 3159 369
rect 3193 335 3199 369
rect 3153 297 3199 335
rect 2821 263 2827 297
rect 2781 251 2827 263
rect 3153 263 3159 297
rect 3193 263 3199 297
rect 3153 251 3199 263
rect 632 200 644 234
rect 678 200 780 234
rect 814 200 826 234
rect 632 194 826 200
rect 548 101 554 135
rect 588 101 594 135
rect 548 89 594 101
rect 161 42 207 80
rect 161 8 167 42
rect 201 8 207 42
rect 161 -4 207 8
<< via1 >>
rect 85 297 137 349
rect 149 320 167 349
rect 167 320 201 349
rect 149 297 201 320
rect 336 828 388 872
rect 336 820 370 828
rect 370 820 388 828
rect 400 820 452 872
rect 3053 820 3105 872
rect 3117 820 3169 872
rect 3009 409 3021 419
rect 3021 409 3055 419
rect 3055 409 3061 419
rect 638 297 690 349
rect 703 297 755 349
rect 768 297 820 349
rect 3009 367 3061 409
rect 2787 335 2821 349
rect 2821 335 2839 349
rect 2787 297 2839 335
rect 2851 297 2903 349
rect 3009 303 3061 355
<< metal2 >>
rect 330 820 336 872
rect 388 820 400 872
rect 452 820 3053 872
rect 3105 820 3117 872
rect 3169 820 3175 872
rect 3009 419 3061 425
tri 2999 367 3009 377 se
tri 2987 355 2999 367 se
rect 2999 355 3061 367
tri 2981 349 2987 355 se
rect 2987 349 3009 355
rect 79 297 85 349
rect 137 297 149 349
rect 201 297 638 349
rect 690 297 703 349
rect 755 297 768 349
rect 820 297 2787 349
rect 2839 297 2851 349
rect 2903 303 3009 349
rect 2903 297 3061 303
use sky130_fd_pr__nfet_01v8__example_55959141808496  sky130_fd_pr__nfet_01v8__example_55959141808496_0
timestamp 1686671242
transform 0 -1 280 1 0 1034
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808497  sky130_fd_pr__nfet_01v8__example_55959141808497_0
timestamp 1686671242
transform 0 1 80 1 0 1627
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808502  sky130_fd_pr__nfet_01v8__example_55959141808502_0
timestamp 1686671242
transform 0 1 80 1 0 2294
box -1 0 289 1
use sky130_fd_pr__nfet_01v8__example_55959141808503  sky130_fd_pr__nfet_01v8__example_55959141808503_0
timestamp 1686671242
transform 0 1 636 1 0 89
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808503  sky130_fd_pr__nfet_01v8__example_55959141808503_1
timestamp 1686671242
transform 0 1 98 1 0 89
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808503  sky130_fd_pr__nfet_01v8__example_55959141808503_2
timestamp 1686671242
transform 0 1 98 1 0 526
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808500  sky130_fd_pr__pfet_01v8__example_55959141808500_0
timestamp 1686671242
transform 1 0 2832 0 1 250
box -1 0 297 1
<< properties >>
string GDS_END 48495682
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48481370
<< end >>
