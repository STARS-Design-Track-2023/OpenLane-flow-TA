magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< metal3 >>
rect 198 6606 3800 6640
rect 198 6016 218 6606
rect 3748 6016 3800 6606
rect 198 4418 3800 6016
rect 198 3616 256 4418
rect 3754 3616 3800 4418
rect 198 3576 3800 3616
<< via3 >>
rect 218 6016 3748 6606
rect 256 3616 3754 4418
<< metal4 >>
rect 0 13600 4000 18593
rect 0 12410 4000 13300
rect 0 11240 4000 12130
rect 0 10874 4000 10940
rect 0 10218 4000 10814
rect 0 9266 4000 9862
rect 0 9140 4000 9206
rect 0 7910 4000 8840
rect 0 6940 4000 7630
rect 0 6606 4000 6660
rect 0 6016 218 6606
rect 3748 6016 4000 6606
rect 0 5970 4000 6016
rect 0 4760 4000 5690
rect 0 4418 4000 4480
rect 0 3616 256 4418
rect 3754 3616 4000 4418
rect 0 3550 4000 3616
rect 0 2580 4000 3270
rect 0 1370 4000 2300
rect 0 0 4000 1090
<< obsm4 >>
rect 0 34750 4000 39593
rect 0 9922 4000 10158
<< metal5 >>
rect 0 34750 4000 39593
rect 0 13600 4000 18590
rect 0 12430 4000 13280
rect 0 11260 4000 12110
rect 0 9140 4000 10940
rect 0 7930 4000 8820
rect 0 6960 4000 7610
rect 0 5990 4000 6640
rect 0 4780 4000 5670
rect 0 3570 4000 4460
rect 0 2600 4000 3250
rect 0 20 4000 2280
<< labels >>
rlabel metal4 s 0 10218 4000 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9266 4000 9862 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 0 9140 4000 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10874 4000 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9140 4000 9206 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6960 4000 7610 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 6940 4000 7630 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 2600 4000 3250 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 2580 4000 3270 6 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 0 5990 4000 6640 6 VSWITCH
port 17 nsew power bidirectional
rlabel metal4 s 0 3550 4000 4480 6 VSWITCH
port 17 nsew power bidirectional
rlabel metal4 s 0 5970 4000 6660 6 VSWITCH
port 17 nsew power bidirectional
rlabel via3 s 256 3616 3754 4418 6 VSWITCH
port 17 nsew power bidirectional
rlabel via3 s 218 6016 3748 6606 6 VSWITCH
port 17 nsew power bidirectional
rlabel metal3 s 198 3576 3800 6640 6 VSWITCH
port 17 nsew power bidirectional
rlabel metal5 s 0 12430 4000 13280 6 VDDIO_Q
port 5 nsew power bidirectional
rlabel metal4 s 0 12410 4000 13300 6 VDDIO_Q
port 5 nsew power bidirectional
rlabel metal5 s 0 20 4000 2280 6 VCCHIB
port 19 nsew power bidirectional
rlabel metal4 s 0 0 4000 1090 6 VCCHIB
port 19 nsew power bidirectional
rlabel metal5 s 0 13600 4000 18590 6 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 0 13600 4000 18593 6 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 0 3570 4000 4460 6 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 0 1370 4000 2300 6 VCCD
port 7 nsew power bidirectional
rlabel metal5 s 0 4780 4000 5670 6 VSSIO
port 8 nsew ground bidirectional
rlabel metal4 s 0 4760 4000 5690 6 VSSIO
port 8 nsew ground bidirectional
rlabel metal5 s 0 34750 4000 39593 6 VSSIO
port 8 nsew ground bidirectional
rlabel metal5 s 0 7930 4000 8820 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 0 7910 4000 8840 6 VSSD
port 9 nsew ground bidirectional
rlabel metal5 s 0 11260 4000 12110 6 VSSIO_Q
port 10 nsew ground bidirectional
rlabel metal4 s 0 11240 4000 12130 6 VSSIO_Q
port 10 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 4000 39593
string LEFclass PAD AREAIO
string LEFview TRUE
string GDS_END 56710
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um.gds
string GDS_START 214
<< end >>
