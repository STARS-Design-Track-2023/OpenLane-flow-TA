magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< locali >>
rect 181 1140 189 1174
rect 223 1140 261 1174
rect 295 1140 333 1174
rect 367 1140 405 1174
rect 439 1140 477 1174
rect 511 1140 519 1174
rect 181 20 189 54
rect 223 20 261 54
rect 295 20 333 54
rect 367 20 405 54
rect 439 20 477 54
rect 511 20 519 54
<< viali >>
rect 189 1140 223 1174
rect 261 1140 295 1174
rect 333 1140 367 1174
rect 405 1140 439 1174
rect 477 1140 511 1174
rect 189 20 223 54
rect 261 20 295 54
rect 333 20 367 54
rect 405 20 439 54
rect 477 20 511 54
<< obsli1 >>
rect 38 1010 72 1048
rect 38 938 72 976
rect 38 866 72 904
rect 38 794 72 832
rect 38 722 72 760
rect 38 650 72 688
rect 38 578 72 616
rect 38 506 72 544
rect 38 434 72 472
rect 38 362 72 400
rect 38 290 72 328
rect 38 218 72 256
rect 38 112 72 184
rect 149 88 183 1106
rect 241 88 275 1106
rect 333 88 367 1106
rect 425 88 459 1106
rect 517 88 551 1106
rect 628 1010 662 1048
rect 628 938 662 976
rect 628 866 662 904
rect 628 794 662 832
rect 628 722 662 760
rect 628 650 662 688
rect 628 578 662 616
rect 628 506 662 544
rect 628 434 662 472
rect 628 362 662 400
rect 628 290 662 328
rect 628 218 662 256
rect 628 112 662 184
<< obsli1c >>
rect 38 1048 72 1082
rect 38 976 72 1010
rect 38 904 72 938
rect 38 832 72 866
rect 38 760 72 794
rect 38 688 72 722
rect 38 616 72 650
rect 38 544 72 578
rect 38 472 72 506
rect 38 400 72 434
rect 38 328 72 362
rect 38 256 72 290
rect 38 184 72 218
rect 628 1048 662 1082
rect 628 976 662 1010
rect 628 904 662 938
rect 628 832 662 866
rect 628 760 662 794
rect 628 688 662 722
rect 628 616 662 650
rect 628 544 662 578
rect 628 472 662 506
rect 628 400 662 434
rect 628 328 662 362
rect 628 256 662 290
rect 628 184 662 218
<< metal1 >>
rect 177 1174 523 1194
rect 177 1140 189 1174
rect 223 1140 261 1174
rect 295 1140 333 1174
rect 367 1140 405 1174
rect 439 1140 477 1174
rect 511 1140 523 1174
rect 177 1128 523 1140
rect 26 1082 84 1094
rect 26 1048 38 1082
rect 72 1048 84 1082
rect 26 1010 84 1048
rect 26 976 38 1010
rect 72 976 84 1010
rect 26 938 84 976
rect 26 904 38 938
rect 72 904 84 938
rect 26 866 84 904
rect 26 832 38 866
rect 72 832 84 866
rect 26 794 84 832
rect 26 760 38 794
rect 72 760 84 794
rect 26 722 84 760
rect 26 688 38 722
rect 72 688 84 722
rect 26 650 84 688
rect 26 616 38 650
rect 72 616 84 650
rect 26 578 84 616
rect 26 544 38 578
rect 72 544 84 578
rect 26 506 84 544
rect 26 472 38 506
rect 72 472 84 506
rect 26 434 84 472
rect 26 400 38 434
rect 72 400 84 434
rect 26 362 84 400
rect 26 328 38 362
rect 72 328 84 362
rect 26 290 84 328
rect 26 256 38 290
rect 72 256 84 290
rect 26 218 84 256
rect 26 184 38 218
rect 72 184 84 218
rect 26 100 84 184
rect 616 1082 674 1094
rect 616 1048 628 1082
rect 662 1048 674 1082
rect 616 1010 674 1048
rect 616 976 628 1010
rect 662 976 674 1010
rect 616 938 674 976
rect 616 904 628 938
rect 662 904 674 938
rect 616 866 674 904
rect 616 832 628 866
rect 662 832 674 866
rect 616 794 674 832
rect 616 760 628 794
rect 662 760 674 794
rect 616 722 674 760
rect 616 688 628 722
rect 662 688 674 722
rect 616 650 674 688
rect 616 616 628 650
rect 662 616 674 650
rect 616 578 674 616
rect 616 544 628 578
rect 662 544 674 578
rect 616 506 674 544
rect 616 472 628 506
rect 662 472 674 506
rect 616 434 674 472
rect 616 400 628 434
rect 662 400 674 434
rect 616 362 674 400
rect 616 328 628 362
rect 662 328 674 362
rect 616 290 674 328
rect 616 256 628 290
rect 662 256 674 290
rect 616 218 674 256
rect 616 184 628 218
rect 662 184 674 218
rect 616 100 674 184
rect 177 54 523 66
rect 177 20 189 54
rect 223 20 261 54
rect 295 20 333 54
rect 367 20 405 54
rect 439 20 477 54
rect 511 20 523 54
rect 177 0 523 20
<< obsm1 >>
rect 140 100 192 1094
rect 232 100 284 1094
rect 324 100 376 1094
rect 416 100 468 1094
rect 508 100 560 1094
<< metal2 >>
rect 0 622 700 1094
rect 0 100 700 572
<< labels >>
rlabel metal2 s 0 622 700 1094 6 DRAIN
port 1 nsew
rlabel viali s 477 1140 511 1174 6 GATE
port 2 nsew
rlabel viali s 477 20 511 54 6 GATE
port 2 nsew
rlabel viali s 405 1140 439 1174 6 GATE
port 2 nsew
rlabel viali s 405 20 439 54 6 GATE
port 2 nsew
rlabel viali s 333 1140 367 1174 6 GATE
port 2 nsew
rlabel viali s 333 20 367 54 6 GATE
port 2 nsew
rlabel viali s 261 1140 295 1174 6 GATE
port 2 nsew
rlabel viali s 261 20 295 54 6 GATE
port 2 nsew
rlabel viali s 189 1140 223 1174 6 GATE
port 2 nsew
rlabel viali s 189 20 223 54 6 GATE
port 2 nsew
rlabel locali s 181 1140 519 1174 6 GATE
port 2 nsew
rlabel locali s 181 20 519 54 6 GATE
port 2 nsew
rlabel metal1 s 177 1128 523 1194 6 GATE
port 2 nsew
rlabel metal1 s 177 0 523 66 6 GATE
port 2 nsew
rlabel metal2 s 0 100 700 572 6 SOURCE
port 3 nsew
rlabel metal1 s 26 100 84 1094 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 616 100 674 1094 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 700 1194
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6116650
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6094560
<< end >>
