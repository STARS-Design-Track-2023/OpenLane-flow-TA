magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1195 203
rect 30 -17 64 21
<< locali >>
rect 103 391 169 425
rect 119 325 153 391
rect 287 325 321 425
rect 29 257 65 325
rect 119 291 436 325
rect 29 215 165 257
rect 209 216 345 257
rect 235 215 301 216
rect 393 165 436 291
rect 483 215 644 325
rect 745 215 896 325
rect 943 215 1172 325
rect 271 131 620 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 35 459 405 493
rect 35 359 69 459
rect 203 359 237 459
rect 371 417 405 459
rect 454 451 588 527
rect 636 417 670 493
rect 710 451 844 527
rect 878 417 912 493
rect 953 451 1087 527
rect 1127 417 1161 493
rect 371 383 1161 417
rect 371 359 405 383
rect 636 359 670 383
rect 878 359 912 383
rect 1127 359 1161 383
rect 35 143 237 177
rect 35 93 69 143
rect 19 59 85 93
rect 119 17 153 109
rect 203 93 237 143
rect 724 127 1078 161
rect 187 59 423 93
rect 470 59 874 93
rect 911 17 978 93
rect 1012 55 1078 127
rect 1112 17 1177 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 483 215 644 325 6 A1
port 1 nsew signal input
rlabel locali s 745 215 896 325 6 A2
port 2 nsew signal input
rlabel locali s 943 215 1172 325 6 A3
port 3 nsew signal input
rlabel locali s 235 215 301 216 6 B1
port 4 nsew signal input
rlabel locali s 209 216 345 257 6 B1
port 4 nsew signal input
rlabel locali s 29 215 165 257 6 B2
port 5 nsew signal input
rlabel locali s 29 257 65 325 6 B2
port 5 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 1195 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 271 131 620 165 6 Y
port 10 nsew signal output
rlabel locali s 393 165 436 291 6 Y
port 10 nsew signal output
rlabel locali s 119 291 436 325 6 Y
port 10 nsew signal output
rlabel locali s 287 325 321 425 6 Y
port 10 nsew signal output
rlabel locali s 119 325 153 391 6 Y
port 10 nsew signal output
rlabel locali s 103 391 169 425 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3504422
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3493188
<< end >>
