magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__dfl1sd__example_55959141808340  sky130_fd_pr__dfl1sd__example_55959141808340_0
timestamp 1686671242
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808341  sky130_fd_pr__hvdfl1sd2__example_55959141808341_0
timestamp 1686671242
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808341  sky130_fd_pr__hvdfl1sd2__example_55959141808341_1
timestamp 1686671242
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808341  sky130_fd_pr__hvdfl1sd2__example_55959141808341_2
timestamp 1686671242
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808342  sky130_fd_pr__hvdfl1sd__example_55959141808342_0
timestamp 1686671242
transform 1 0 568 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 36943866
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 36941260
<< end >>
