magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 1989 203
rect 27 -17 61 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 419 47 449 177
rect 503 47 533 177
rect 587 47 617 177
rect 671 47 701 177
rect 859 47 889 177
rect 943 47 973 177
rect 1027 47 1057 177
rect 1111 47 1141 177
rect 1293 47 1323 177
rect 1377 47 1407 177
rect 1461 47 1491 177
rect 1545 47 1575 177
rect 1629 47 1659 177
rect 1713 47 1743 177
rect 1797 47 1827 177
rect 1881 47 1911 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 419 297 449 497
rect 503 297 533 497
rect 587 297 617 497
rect 671 297 701 497
rect 853 297 883 497
rect 937 297 967 497
rect 1021 297 1051 497
rect 1105 297 1135 497
rect 1293 297 1323 497
rect 1377 297 1407 497
rect 1461 297 1491 497
rect 1545 297 1575 497
rect 1629 297 1659 497
rect 1713 297 1743 497
rect 1797 297 1827 497
rect 1881 297 1911 497
<< ndiff >>
rect 27 95 83 177
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 47 167 129
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 47 335 129
rect 365 163 419 177
rect 365 129 375 163
rect 409 129 419 163
rect 365 95 419 129
rect 365 61 375 95
rect 409 61 419 95
rect 365 47 419 61
rect 449 95 503 177
rect 449 61 459 95
rect 493 61 503 95
rect 449 47 503 61
rect 533 163 587 177
rect 533 129 543 163
rect 577 129 587 163
rect 533 95 587 129
rect 533 61 543 95
rect 577 61 587 95
rect 533 47 587 61
rect 617 95 671 177
rect 617 61 627 95
rect 661 61 671 95
rect 617 47 671 61
rect 701 163 753 177
rect 701 129 711 163
rect 745 129 753 163
rect 701 95 753 129
rect 701 61 711 95
rect 745 61 753 95
rect 701 47 753 61
rect 807 133 859 177
rect 807 99 815 133
rect 849 99 859 133
rect 807 47 859 99
rect 889 163 943 177
rect 889 129 899 163
rect 933 129 943 163
rect 889 47 943 129
rect 973 95 1027 177
rect 973 61 983 95
rect 1017 61 1027 95
rect 973 47 1027 61
rect 1057 163 1111 177
rect 1057 129 1067 163
rect 1101 129 1111 163
rect 1057 47 1111 129
rect 1141 95 1293 177
rect 1141 61 1151 95
rect 1185 61 1249 95
rect 1283 61 1293 95
rect 1141 47 1293 61
rect 1323 95 1377 177
rect 1323 61 1333 95
rect 1367 61 1377 95
rect 1323 47 1377 61
rect 1407 163 1461 177
rect 1407 129 1417 163
rect 1451 129 1461 163
rect 1407 95 1461 129
rect 1407 61 1417 95
rect 1451 61 1461 95
rect 1407 47 1461 61
rect 1491 95 1545 177
rect 1491 61 1501 95
rect 1535 61 1545 95
rect 1491 47 1545 61
rect 1575 163 1629 177
rect 1575 129 1585 163
rect 1619 129 1629 163
rect 1575 95 1629 129
rect 1575 61 1585 95
rect 1619 61 1629 95
rect 1575 47 1629 61
rect 1659 95 1713 177
rect 1659 61 1669 95
rect 1703 61 1713 95
rect 1659 47 1713 61
rect 1743 163 1797 177
rect 1743 129 1753 163
rect 1787 129 1797 163
rect 1743 95 1797 129
rect 1743 61 1753 95
rect 1787 61 1797 95
rect 1743 47 1797 61
rect 1827 95 1881 177
rect 1827 61 1837 95
rect 1871 61 1881 95
rect 1827 47 1881 61
rect 1911 163 1963 177
rect 1911 129 1921 163
rect 1955 129 1963 163
rect 1911 95 1963 129
rect 1911 61 1921 95
rect 1955 61 1963 95
rect 1911 47 1963 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 297 83 375
rect 113 477 167 497
rect 113 443 123 477
rect 157 443 167 477
rect 113 409 167 443
rect 113 375 123 409
rect 157 375 167 409
rect 113 341 167 375
rect 113 307 123 341
rect 157 307 167 341
rect 113 297 167 307
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 297 251 375
rect 281 477 335 497
rect 281 443 291 477
rect 325 443 335 477
rect 281 409 335 443
rect 281 375 291 409
rect 325 375 335 409
rect 281 341 335 375
rect 281 307 291 341
rect 325 307 335 341
rect 281 297 335 307
rect 365 477 419 497
rect 365 443 375 477
rect 409 443 419 477
rect 365 409 419 443
rect 365 375 375 409
rect 409 375 419 409
rect 365 297 419 375
rect 449 477 503 497
rect 449 443 459 477
rect 493 443 503 477
rect 449 409 503 443
rect 449 375 459 409
rect 493 375 503 409
rect 449 341 503 375
rect 449 307 459 341
rect 493 307 503 341
rect 449 297 503 307
rect 533 477 587 497
rect 533 443 543 477
rect 577 443 587 477
rect 533 409 587 443
rect 533 375 543 409
rect 577 375 587 409
rect 533 297 587 375
rect 617 477 671 497
rect 617 443 627 477
rect 661 443 671 477
rect 617 409 671 443
rect 617 375 627 409
rect 661 375 671 409
rect 617 341 671 375
rect 617 307 627 341
rect 661 307 671 341
rect 617 297 671 307
rect 701 477 853 497
rect 701 443 711 477
rect 745 443 809 477
rect 843 443 853 477
rect 701 409 853 443
rect 701 375 711 409
rect 745 375 809 409
rect 843 375 853 409
rect 701 297 853 375
rect 883 477 937 497
rect 883 443 893 477
rect 927 443 937 477
rect 883 409 937 443
rect 883 375 893 409
rect 927 375 937 409
rect 883 341 937 375
rect 883 307 893 341
rect 927 307 937 341
rect 883 297 937 307
rect 967 477 1021 497
rect 967 443 977 477
rect 1011 443 1021 477
rect 967 409 1021 443
rect 967 375 977 409
rect 1011 375 1021 409
rect 967 297 1021 375
rect 1051 477 1105 497
rect 1051 443 1061 477
rect 1095 443 1105 477
rect 1051 409 1105 443
rect 1051 375 1061 409
rect 1095 375 1105 409
rect 1051 341 1105 375
rect 1051 307 1061 341
rect 1095 307 1105 341
rect 1051 297 1105 307
rect 1135 477 1187 497
rect 1135 443 1145 477
rect 1179 443 1187 477
rect 1135 409 1187 443
rect 1135 375 1145 409
rect 1179 375 1187 409
rect 1135 297 1187 375
rect 1241 477 1293 497
rect 1241 443 1249 477
rect 1283 443 1293 477
rect 1241 409 1293 443
rect 1241 375 1249 409
rect 1283 375 1293 409
rect 1241 297 1293 375
rect 1323 409 1377 497
rect 1323 375 1333 409
rect 1367 375 1377 409
rect 1323 341 1377 375
rect 1323 307 1333 341
rect 1367 307 1377 341
rect 1323 297 1377 307
rect 1407 477 1461 497
rect 1407 443 1417 477
rect 1451 443 1461 477
rect 1407 409 1461 443
rect 1407 375 1417 409
rect 1451 375 1461 409
rect 1407 297 1461 375
rect 1491 409 1545 497
rect 1491 375 1501 409
rect 1535 375 1545 409
rect 1491 341 1545 375
rect 1491 307 1501 341
rect 1535 307 1545 341
rect 1491 297 1545 307
rect 1575 477 1629 497
rect 1575 443 1585 477
rect 1619 443 1629 477
rect 1575 409 1629 443
rect 1575 375 1585 409
rect 1619 375 1629 409
rect 1575 341 1629 375
rect 1575 307 1585 341
rect 1619 307 1629 341
rect 1575 297 1629 307
rect 1659 477 1713 497
rect 1659 443 1669 477
rect 1703 443 1713 477
rect 1659 409 1713 443
rect 1659 375 1669 409
rect 1703 375 1713 409
rect 1659 297 1713 375
rect 1743 477 1797 497
rect 1743 443 1753 477
rect 1787 443 1797 477
rect 1743 409 1797 443
rect 1743 375 1753 409
rect 1787 375 1797 409
rect 1743 341 1797 375
rect 1743 307 1753 341
rect 1787 307 1797 341
rect 1743 297 1797 307
rect 1827 477 1881 497
rect 1827 443 1837 477
rect 1871 443 1881 477
rect 1827 409 1881 443
rect 1827 375 1837 409
rect 1871 375 1881 409
rect 1827 297 1881 375
rect 1911 477 1967 497
rect 1911 443 1921 477
rect 1955 443 1967 477
rect 1911 409 1967 443
rect 1911 375 1921 409
rect 1955 375 1967 409
rect 1911 341 1967 375
rect 1911 307 1921 341
rect 1955 307 1967 341
rect 1911 297 1967 307
<< ndiffc >>
rect 39 61 73 95
rect 123 129 157 163
rect 207 61 241 95
rect 291 129 325 163
rect 375 129 409 163
rect 375 61 409 95
rect 459 61 493 95
rect 543 129 577 163
rect 543 61 577 95
rect 627 61 661 95
rect 711 129 745 163
rect 711 61 745 95
rect 815 99 849 133
rect 899 129 933 163
rect 983 61 1017 95
rect 1067 129 1101 163
rect 1151 61 1185 95
rect 1249 61 1283 95
rect 1333 61 1367 95
rect 1417 129 1451 163
rect 1417 61 1451 95
rect 1501 61 1535 95
rect 1585 129 1619 163
rect 1585 61 1619 95
rect 1669 61 1703 95
rect 1753 129 1787 163
rect 1753 61 1787 95
rect 1837 61 1871 95
rect 1921 129 1955 163
rect 1921 61 1955 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 123 443 157 477
rect 123 375 157 409
rect 123 307 157 341
rect 207 443 241 477
rect 207 375 241 409
rect 291 443 325 477
rect 291 375 325 409
rect 291 307 325 341
rect 375 443 409 477
rect 375 375 409 409
rect 459 443 493 477
rect 459 375 493 409
rect 459 307 493 341
rect 543 443 577 477
rect 543 375 577 409
rect 627 443 661 477
rect 627 375 661 409
rect 627 307 661 341
rect 711 443 745 477
rect 809 443 843 477
rect 711 375 745 409
rect 809 375 843 409
rect 893 443 927 477
rect 893 375 927 409
rect 893 307 927 341
rect 977 443 1011 477
rect 977 375 1011 409
rect 1061 443 1095 477
rect 1061 375 1095 409
rect 1061 307 1095 341
rect 1145 443 1179 477
rect 1145 375 1179 409
rect 1249 443 1283 477
rect 1249 375 1283 409
rect 1333 375 1367 409
rect 1333 307 1367 341
rect 1417 443 1451 477
rect 1417 375 1451 409
rect 1501 375 1535 409
rect 1501 307 1535 341
rect 1585 443 1619 477
rect 1585 375 1619 409
rect 1585 307 1619 341
rect 1669 443 1703 477
rect 1669 375 1703 409
rect 1753 443 1787 477
rect 1753 375 1787 409
rect 1753 307 1787 341
rect 1837 443 1871 477
rect 1837 375 1871 409
rect 1921 443 1955 477
rect 1921 375 1955 409
rect 1921 307 1955 341
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 419 497 449 523
rect 503 497 533 523
rect 587 497 617 523
rect 671 497 701 523
rect 853 497 883 523
rect 937 497 967 523
rect 1021 497 1051 523
rect 1105 497 1135 523
rect 1293 497 1323 523
rect 1377 497 1407 523
rect 1461 497 1491 523
rect 1545 497 1575 523
rect 1629 497 1659 523
rect 1713 497 1743 523
rect 1797 497 1827 523
rect 1881 497 1911 523
rect 83 265 113 297
rect 167 265 197 297
rect 251 265 281 297
rect 335 265 365 297
rect 83 249 365 265
rect 83 215 101 249
rect 135 215 169 249
rect 203 215 237 249
rect 271 215 305 249
rect 339 215 365 249
rect 83 199 365 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 177 281 199
rect 335 177 365 199
rect 419 265 449 297
rect 503 265 533 297
rect 587 265 617 297
rect 671 265 701 297
rect 419 249 701 265
rect 419 215 435 249
rect 469 215 503 249
rect 537 215 571 249
rect 605 215 639 249
rect 673 215 701 249
rect 419 199 701 215
rect 853 265 883 297
rect 937 265 967 297
rect 1021 265 1051 297
rect 1105 265 1135 297
rect 1293 265 1323 297
rect 1377 265 1407 297
rect 1461 265 1491 297
rect 1545 265 1575 297
rect 853 249 1141 265
rect 853 215 875 249
rect 909 215 943 249
rect 977 215 1011 249
rect 1045 215 1079 249
rect 1113 215 1141 249
rect 853 199 1141 215
rect 419 177 449 199
rect 503 177 533 199
rect 587 177 617 199
rect 671 177 701 199
rect 859 177 889 199
rect 943 177 973 199
rect 1027 177 1057 199
rect 1111 177 1141 199
rect 1293 249 1575 265
rect 1293 215 1309 249
rect 1343 215 1377 249
rect 1411 215 1445 249
rect 1479 215 1513 249
rect 1547 215 1575 249
rect 1293 199 1575 215
rect 1293 177 1323 199
rect 1377 177 1407 199
rect 1461 177 1491 199
rect 1545 177 1575 199
rect 1629 265 1659 297
rect 1713 265 1743 297
rect 1797 265 1827 297
rect 1881 265 1911 297
rect 1629 249 1911 265
rect 1629 215 1639 249
rect 1673 215 1707 249
rect 1741 215 1775 249
rect 1809 215 1843 249
rect 1877 215 1911 249
rect 1629 199 1911 215
rect 1629 177 1659 199
rect 1713 177 1743 199
rect 1797 177 1827 199
rect 1881 177 1911 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 419 21 449 47
rect 503 21 533 47
rect 587 21 617 47
rect 671 21 701 47
rect 859 21 889 47
rect 943 21 973 47
rect 1027 21 1057 47
rect 1111 21 1141 47
rect 1293 21 1323 47
rect 1377 21 1407 47
rect 1461 21 1491 47
rect 1545 21 1575 47
rect 1629 21 1659 47
rect 1713 21 1743 47
rect 1797 21 1827 47
rect 1881 21 1911 47
<< polycont >>
rect 101 215 135 249
rect 169 215 203 249
rect 237 215 271 249
rect 305 215 339 249
rect 435 215 469 249
rect 503 215 537 249
rect 571 215 605 249
rect 639 215 673 249
rect 875 215 909 249
rect 943 215 977 249
rect 1011 215 1045 249
rect 1079 215 1113 249
rect 1309 215 1343 249
rect 1377 215 1411 249
rect 1445 215 1479 249
rect 1513 215 1547 249
rect 1639 215 1673 249
rect 1707 215 1741 249
rect 1775 215 1809 249
rect 1843 215 1877 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 31 477 81 527
rect 31 443 39 477
rect 73 443 81 477
rect 31 409 81 443
rect 31 375 39 409
rect 73 375 81 409
rect 31 359 81 375
rect 115 477 165 493
rect 115 443 123 477
rect 157 443 165 477
rect 115 409 165 443
rect 115 375 123 409
rect 157 375 165 409
rect 115 341 165 375
rect 199 477 249 527
rect 199 443 207 477
rect 241 443 249 477
rect 199 409 249 443
rect 199 375 207 409
rect 241 375 249 409
rect 199 359 249 375
rect 283 477 333 493
rect 283 443 291 477
rect 325 443 333 477
rect 283 409 333 443
rect 283 375 291 409
rect 325 375 333 409
rect 115 325 123 341
rect 17 307 123 325
rect 157 325 165 341
rect 283 341 333 375
rect 367 477 417 527
rect 367 443 375 477
rect 409 443 417 477
rect 367 409 417 443
rect 367 375 375 409
rect 409 375 417 409
rect 367 359 417 375
rect 451 477 501 493
rect 451 443 459 477
rect 493 443 501 477
rect 451 409 501 443
rect 451 375 459 409
rect 493 375 501 409
rect 283 325 291 341
rect 157 307 291 325
rect 325 325 333 341
rect 451 341 501 375
rect 535 477 585 527
rect 535 443 543 477
rect 577 443 585 477
rect 535 409 585 443
rect 535 375 543 409
rect 577 375 585 409
rect 535 359 585 375
rect 619 477 669 493
rect 619 443 627 477
rect 661 443 669 477
rect 619 409 669 443
rect 619 375 627 409
rect 661 375 669 409
rect 451 325 459 341
rect 325 307 459 325
rect 493 325 501 341
rect 619 341 669 375
rect 703 477 851 527
rect 703 443 711 477
rect 745 443 809 477
rect 843 443 851 477
rect 703 409 851 443
rect 703 375 711 409
rect 745 375 809 409
rect 843 375 851 409
rect 703 359 851 375
rect 885 477 935 493
rect 885 443 893 477
rect 927 443 935 477
rect 885 409 935 443
rect 885 375 893 409
rect 927 375 935 409
rect 619 325 627 341
rect 493 307 627 325
rect 661 325 669 341
rect 885 341 935 375
rect 969 477 1019 527
rect 969 443 977 477
rect 1011 443 1019 477
rect 969 409 1019 443
rect 969 375 977 409
rect 1011 375 1019 409
rect 969 359 1019 375
rect 1053 477 1103 493
rect 1053 443 1061 477
rect 1095 443 1103 477
rect 1053 409 1103 443
rect 1053 375 1061 409
rect 1095 375 1103 409
rect 661 307 783 325
rect 17 291 783 307
rect 885 307 893 341
rect 927 325 935 341
rect 1053 341 1103 375
rect 1137 477 1187 527
rect 1137 443 1145 477
rect 1179 443 1187 477
rect 1137 409 1187 443
rect 1137 375 1145 409
rect 1179 375 1187 409
rect 1137 359 1187 375
rect 1235 477 1627 493
rect 1235 443 1249 477
rect 1283 459 1417 477
rect 1283 443 1291 459
rect 1235 409 1291 443
rect 1409 443 1417 459
rect 1451 459 1585 477
rect 1451 443 1459 459
rect 1235 375 1249 409
rect 1283 375 1291 409
rect 1235 359 1291 375
rect 1325 409 1375 425
rect 1325 375 1333 409
rect 1367 375 1375 409
rect 1053 325 1061 341
rect 927 307 1061 325
rect 1095 325 1103 341
rect 1325 341 1375 375
rect 1409 409 1459 443
rect 1577 443 1585 459
rect 1619 443 1627 477
rect 1409 375 1417 409
rect 1451 375 1459 409
rect 1409 359 1459 375
rect 1493 409 1543 425
rect 1493 375 1501 409
rect 1535 375 1543 409
rect 1325 325 1333 341
rect 1095 307 1333 325
rect 1367 325 1375 341
rect 1493 341 1543 375
rect 1493 325 1501 341
rect 1367 307 1501 325
rect 1535 307 1543 341
rect 885 291 1543 307
rect 1577 409 1627 443
rect 1577 375 1585 409
rect 1619 375 1627 409
rect 1577 341 1627 375
rect 1661 477 1711 527
rect 1661 443 1669 477
rect 1703 443 1711 477
rect 1661 409 1711 443
rect 1661 375 1669 409
rect 1703 375 1711 409
rect 1661 359 1711 375
rect 1745 477 1795 493
rect 1745 443 1753 477
rect 1787 443 1795 477
rect 1745 409 1795 443
rect 1745 375 1753 409
rect 1787 375 1795 409
rect 1577 307 1585 341
rect 1619 325 1627 341
rect 1745 341 1795 375
rect 1829 477 1879 527
rect 1829 443 1837 477
rect 1871 443 1879 477
rect 1829 409 1879 443
rect 1829 375 1837 409
rect 1871 375 1879 409
rect 1829 359 1879 375
rect 1913 477 1975 493
rect 1913 443 1921 477
rect 1955 443 1975 477
rect 1913 409 1975 443
rect 1913 375 1921 409
rect 1955 375 1975 409
rect 1745 325 1753 341
rect 1619 307 1753 325
rect 1787 325 1795 341
rect 1913 341 1975 375
rect 1913 325 1921 341
rect 1787 307 1921 325
rect 1955 307 1975 341
rect 1577 291 1975 307
rect 17 181 51 291
rect 749 257 783 291
rect 85 249 365 257
rect 85 215 101 249
rect 135 215 169 249
rect 203 215 237 249
rect 271 215 305 249
rect 339 215 365 249
rect 419 249 701 257
rect 419 215 435 249
rect 469 215 503 249
rect 537 215 571 249
rect 605 215 639 249
rect 673 215 701 249
rect 749 249 1141 257
rect 749 215 875 249
rect 909 215 943 249
rect 977 215 1011 249
rect 1045 215 1079 249
rect 1113 215 1141 249
rect 1175 181 1231 291
rect 1293 249 1575 257
rect 1293 215 1309 249
rect 1343 215 1377 249
rect 1411 215 1445 249
rect 1479 215 1513 249
rect 1547 215 1575 249
rect 1609 249 2001 257
rect 1609 215 1639 249
rect 1673 215 1707 249
rect 1741 215 1775 249
rect 1809 215 1843 249
rect 1877 215 2001 249
rect 17 163 341 181
rect 17 129 123 163
rect 157 129 291 163
rect 325 129 341 163
rect 375 163 761 181
rect 409 145 543 163
rect 409 129 425 145
rect 375 95 425 129
rect 527 129 543 145
rect 577 145 711 163
rect 577 129 593 145
rect 20 61 39 95
rect 73 61 207 95
rect 241 61 375 95
rect 409 61 425 95
rect 20 51 425 61
rect 459 95 493 111
rect 459 17 493 61
rect 527 95 593 129
rect 695 129 711 145
rect 745 129 761 163
rect 527 61 543 95
rect 577 61 593 95
rect 527 51 593 61
rect 627 95 661 111
rect 627 17 661 61
rect 695 95 761 129
rect 695 61 711 95
rect 745 61 761 95
rect 695 51 761 61
rect 812 133 849 167
rect 812 99 815 133
rect 883 163 1231 181
rect 883 129 899 163
rect 933 129 1067 163
rect 1101 129 1231 163
rect 1265 163 1971 181
rect 1265 147 1417 163
rect 812 95 849 99
rect 1265 95 1299 147
rect 1401 129 1417 147
rect 1451 145 1585 163
rect 1451 129 1467 145
rect 812 61 983 95
rect 1017 61 1151 95
rect 1185 61 1249 95
rect 1283 61 1299 95
rect 812 51 1299 61
rect 1333 95 1367 111
rect 1333 17 1367 61
rect 1401 95 1467 129
rect 1569 129 1585 145
rect 1619 145 1753 163
rect 1619 129 1635 145
rect 1401 61 1417 95
rect 1451 61 1467 95
rect 1401 51 1467 61
rect 1501 95 1535 111
rect 1501 17 1535 61
rect 1569 95 1635 129
rect 1737 129 1753 145
rect 1787 145 1921 163
rect 1787 129 1803 145
rect 1569 61 1585 95
rect 1619 61 1635 95
rect 1569 51 1635 61
rect 1669 95 1703 111
rect 1669 17 1703 61
rect 1737 95 1803 129
rect 1905 129 1921 145
rect 1955 129 1971 163
rect 1737 61 1753 95
rect 1787 61 1803 95
rect 1737 51 1803 61
rect 1837 95 1871 111
rect 1837 17 1871 61
rect 1905 95 1971 129
rect 1905 61 1921 95
rect 1955 61 1971 95
rect 1905 51 1971 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 579 221 613 255 0 FreeSans 400 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 1777 221 1811 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 1409 221 1443 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 211 221 245 255 0 FreeSans 400 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 1501 357 1535 391 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel nwell s 27 527 61 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 27 -17 61 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 27 -17 61 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 27 527 61 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o2bb2ai_4
rlabel metal1 s 0 -48 2024 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2024 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 1264842
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1250080
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 10.120 0.000 
<< end >>
