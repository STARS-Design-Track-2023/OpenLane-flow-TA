magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 5 13 363 203
rect 35 -12 57 13
<< ndiff >>
rect 31 39 337 177
<< pdiff >>
rect 31 305 337 505
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel metal1 s 34 -10 57 9 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 34 535 54 552 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 35 530 60 556 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 35 -12 57 12 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 fill_4
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_END 3954636
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3952896
string path 0.000 0.000 9.200 0.000 
<< end >>
