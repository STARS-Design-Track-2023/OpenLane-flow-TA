magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect 7177 3556 11455 3812
rect 7177 396 7483 3556
rect 11159 396 11455 3556
rect 7177 140 11455 396
<< pwell >>
rect 7497 450 11145 3502
<< mvpsubdiff >>
rect 7523 3421 7823 3476
rect 7523 531 7554 3421
rect 7792 531 7823 3421
rect 7523 476 7823 531
rect 8347 3421 8647 3476
rect 8347 531 8378 3421
rect 8616 531 8647 3421
rect 8347 476 8647 531
rect 9171 3421 9471 3476
rect 9171 531 9202 3421
rect 9440 531 9471 3421
rect 9171 476 9471 531
rect 9995 3421 10295 3476
rect 9995 531 10026 3421
rect 10264 531 10295 3421
rect 9995 476 10295 531
rect 10819 3421 11119 3476
rect 10819 531 10850 3421
rect 11088 531 11119 3421
rect 10819 476 11119 531
<< mvnsubdiff >>
rect 7243 3694 11389 3746
rect 7243 3660 7353 3694
rect 7387 3660 7421 3694
rect 7455 3660 7489 3694
rect 7523 3660 7557 3694
rect 7591 3660 7625 3694
rect 7659 3660 7693 3694
rect 7727 3660 7761 3694
rect 7795 3660 7829 3694
rect 7863 3660 7897 3694
rect 7931 3660 7965 3694
rect 7999 3660 8033 3694
rect 8067 3660 8101 3694
rect 8135 3660 8169 3694
rect 8203 3660 8237 3694
rect 8271 3660 8305 3694
rect 8339 3660 8373 3694
rect 8407 3660 8441 3694
rect 8475 3660 8509 3694
rect 8543 3660 8577 3694
rect 8611 3660 8645 3694
rect 8679 3660 8713 3694
rect 8747 3660 8781 3694
rect 8815 3660 8849 3694
rect 8883 3660 8917 3694
rect 8951 3660 8985 3694
rect 9019 3660 9053 3694
rect 9087 3660 9121 3694
rect 9155 3660 9189 3694
rect 9223 3660 9257 3694
rect 9291 3660 9325 3694
rect 9359 3660 9393 3694
rect 9427 3660 9461 3694
rect 9495 3660 9529 3694
rect 9563 3660 9597 3694
rect 9631 3660 9665 3694
rect 9699 3660 9733 3694
rect 9767 3660 9801 3694
rect 9835 3660 9869 3694
rect 9903 3660 9937 3694
rect 9971 3660 10005 3694
rect 10039 3660 10073 3694
rect 10107 3660 10141 3694
rect 10175 3660 10209 3694
rect 10243 3660 10277 3694
rect 10311 3660 10345 3694
rect 10379 3660 10413 3694
rect 10447 3660 10481 3694
rect 10515 3660 10549 3694
rect 10583 3660 10617 3694
rect 10651 3660 10685 3694
rect 10719 3660 10753 3694
rect 10787 3660 10821 3694
rect 10855 3660 10889 3694
rect 10923 3660 10957 3694
rect 10991 3660 11025 3694
rect 11059 3660 11093 3694
rect 11127 3660 11161 3694
rect 11195 3660 11229 3694
rect 11263 3660 11389 3694
rect 7243 3628 11389 3660
rect 7243 3557 7371 3628
rect 7243 3523 7277 3557
rect 7311 3523 7371 3557
rect 7243 3489 7371 3523
rect 7243 3455 7277 3489
rect 7311 3455 7371 3489
rect 11271 3557 11389 3628
rect 11271 3523 11331 3557
rect 11365 3523 11389 3557
rect 11271 3489 11389 3523
rect 7243 3421 7371 3455
rect 7243 3387 7277 3421
rect 7311 3387 7371 3421
rect 7243 3353 7371 3387
rect 7243 3319 7277 3353
rect 7311 3319 7371 3353
rect 7243 3285 7371 3319
rect 7243 3251 7277 3285
rect 7311 3251 7371 3285
rect 7243 3217 7371 3251
rect 7243 3183 7277 3217
rect 7311 3183 7371 3217
rect 7243 3149 7371 3183
rect 7243 3115 7277 3149
rect 7311 3115 7371 3149
rect 7243 3081 7371 3115
rect 7243 3047 7277 3081
rect 7311 3047 7371 3081
rect 7243 3013 7371 3047
rect 7243 2979 7277 3013
rect 7311 2979 7371 3013
rect 7243 2945 7371 2979
rect 7243 2911 7277 2945
rect 7311 2911 7371 2945
rect 7243 2877 7371 2911
rect 7243 2843 7277 2877
rect 7311 2843 7371 2877
rect 7243 2809 7371 2843
rect 7243 2775 7277 2809
rect 7311 2775 7371 2809
rect 7243 2741 7371 2775
rect 7243 2707 7277 2741
rect 7311 2707 7371 2741
rect 7243 2673 7371 2707
rect 7243 2639 7277 2673
rect 7311 2639 7371 2673
rect 7243 2605 7371 2639
rect 7243 2571 7277 2605
rect 7311 2571 7371 2605
rect 7243 2537 7371 2571
rect 7243 2503 7277 2537
rect 7311 2503 7371 2537
rect 7243 2469 7371 2503
rect 7243 2435 7277 2469
rect 7311 2435 7371 2469
rect 7243 2401 7371 2435
rect 7243 2367 7277 2401
rect 7311 2367 7371 2401
rect 7243 2333 7371 2367
rect 7243 2299 7277 2333
rect 7311 2299 7371 2333
rect 7243 2265 7371 2299
rect 7243 2231 7277 2265
rect 7311 2231 7371 2265
rect 7243 2197 7371 2231
rect 7243 2163 7277 2197
rect 7311 2163 7371 2197
rect 7243 2129 7371 2163
rect 7243 2095 7277 2129
rect 7311 2095 7371 2129
rect 7243 2061 7371 2095
rect 7243 2027 7277 2061
rect 7311 2027 7371 2061
rect 7243 1993 7371 2027
rect 7243 1959 7277 1993
rect 7311 1959 7371 1993
rect 7243 1925 7371 1959
rect 7243 1891 7277 1925
rect 7311 1891 7371 1925
rect 7243 1857 7371 1891
rect 7243 1823 7277 1857
rect 7311 1823 7371 1857
rect 7243 1789 7371 1823
rect 7243 1755 7277 1789
rect 7311 1755 7371 1789
rect 7243 1721 7371 1755
rect 7243 1687 7277 1721
rect 7311 1687 7371 1721
rect 7243 1653 7371 1687
rect 7243 1619 7277 1653
rect 7311 1619 7371 1653
rect 7243 1585 7371 1619
rect 7243 1551 7277 1585
rect 7311 1551 7371 1585
rect 7243 1517 7371 1551
rect 7243 1483 7277 1517
rect 7311 1483 7371 1517
rect 7243 1449 7371 1483
rect 7243 1415 7277 1449
rect 7311 1415 7371 1449
rect 7243 1381 7371 1415
rect 7243 1347 7277 1381
rect 7311 1347 7371 1381
rect 7243 1313 7371 1347
rect 7243 1279 7277 1313
rect 7311 1279 7371 1313
rect 7243 1245 7371 1279
rect 7243 1211 7277 1245
rect 7311 1211 7371 1245
rect 7243 1177 7371 1211
rect 7243 1143 7277 1177
rect 7311 1143 7371 1177
rect 7243 1109 7371 1143
rect 7243 1075 7277 1109
rect 7311 1075 7371 1109
rect 7243 1041 7371 1075
rect 7243 1007 7277 1041
rect 7311 1007 7371 1041
rect 7243 973 7371 1007
rect 7243 939 7277 973
rect 7311 939 7371 973
rect 7243 905 7371 939
rect 7243 871 7277 905
rect 7311 871 7371 905
rect 7243 837 7371 871
rect 7243 803 7277 837
rect 7311 803 7371 837
rect 7243 769 7371 803
rect 7243 735 7277 769
rect 7311 735 7371 769
rect 7243 701 7371 735
rect 7243 667 7277 701
rect 7311 667 7371 701
rect 7243 633 7371 667
rect 7243 599 7277 633
rect 7311 599 7371 633
rect 7243 565 7371 599
rect 7243 531 7277 565
rect 7311 531 7371 565
rect 7243 497 7371 531
rect 7243 463 7277 497
rect 7311 463 7371 497
rect 11271 3455 11331 3489
rect 11365 3455 11389 3489
rect 11271 3421 11389 3455
rect 11271 3387 11331 3421
rect 11365 3387 11389 3421
rect 11271 3353 11389 3387
rect 11271 3319 11331 3353
rect 11365 3319 11389 3353
rect 11271 3285 11389 3319
rect 11271 3251 11331 3285
rect 11365 3251 11389 3285
rect 11271 3217 11389 3251
rect 11271 3183 11331 3217
rect 11365 3183 11389 3217
rect 11271 3149 11389 3183
rect 11271 3115 11331 3149
rect 11365 3115 11389 3149
rect 11271 3081 11389 3115
rect 11271 3047 11331 3081
rect 11365 3047 11389 3081
rect 11271 3013 11389 3047
rect 11271 2979 11331 3013
rect 11365 2979 11389 3013
rect 11271 2945 11389 2979
rect 11271 2911 11331 2945
rect 11365 2911 11389 2945
rect 11271 2877 11389 2911
rect 11271 2843 11331 2877
rect 11365 2843 11389 2877
rect 11271 2809 11389 2843
rect 11271 2775 11331 2809
rect 11365 2775 11389 2809
rect 11271 2741 11389 2775
rect 11271 2707 11331 2741
rect 11365 2707 11389 2741
rect 11271 2673 11389 2707
rect 11271 2639 11331 2673
rect 11365 2639 11389 2673
rect 11271 2605 11389 2639
rect 11271 2571 11331 2605
rect 11365 2571 11389 2605
rect 11271 2537 11389 2571
rect 11271 2503 11331 2537
rect 11365 2503 11389 2537
rect 11271 2469 11389 2503
rect 11271 2435 11331 2469
rect 11365 2435 11389 2469
rect 11271 2401 11389 2435
rect 11271 2367 11331 2401
rect 11365 2367 11389 2401
rect 11271 2333 11389 2367
rect 11271 2299 11331 2333
rect 11365 2299 11389 2333
rect 11271 2265 11389 2299
rect 11271 2231 11331 2265
rect 11365 2231 11389 2265
rect 11271 2197 11389 2231
rect 11271 2163 11331 2197
rect 11365 2163 11389 2197
rect 11271 2129 11389 2163
rect 11271 2095 11331 2129
rect 11365 2095 11389 2129
rect 11271 2061 11389 2095
rect 11271 2027 11331 2061
rect 11365 2027 11389 2061
rect 11271 1993 11389 2027
rect 11271 1959 11331 1993
rect 11365 1959 11389 1993
rect 11271 1925 11389 1959
rect 11271 1891 11331 1925
rect 11365 1891 11389 1925
rect 11271 1857 11389 1891
rect 11271 1823 11331 1857
rect 11365 1823 11389 1857
rect 11271 1789 11389 1823
rect 11271 1755 11331 1789
rect 11365 1755 11389 1789
rect 11271 1721 11389 1755
rect 11271 1687 11331 1721
rect 11365 1687 11389 1721
rect 11271 1653 11389 1687
rect 11271 1619 11331 1653
rect 11365 1619 11389 1653
rect 11271 1585 11389 1619
rect 11271 1551 11331 1585
rect 11365 1551 11389 1585
rect 11271 1517 11389 1551
rect 11271 1483 11331 1517
rect 11365 1483 11389 1517
rect 11271 1449 11389 1483
rect 11271 1415 11331 1449
rect 11365 1415 11389 1449
rect 11271 1381 11389 1415
rect 11271 1347 11331 1381
rect 11365 1347 11389 1381
rect 11271 1313 11389 1347
rect 11271 1279 11331 1313
rect 11365 1279 11389 1313
rect 11271 1245 11389 1279
rect 11271 1211 11331 1245
rect 11365 1211 11389 1245
rect 11271 1177 11389 1211
rect 11271 1143 11331 1177
rect 11365 1143 11389 1177
rect 11271 1109 11389 1143
rect 11271 1075 11331 1109
rect 11365 1075 11389 1109
rect 11271 1041 11389 1075
rect 11271 1007 11331 1041
rect 11365 1007 11389 1041
rect 11271 973 11389 1007
rect 11271 939 11331 973
rect 11365 939 11389 973
rect 11271 905 11389 939
rect 11271 871 11331 905
rect 11365 871 11389 905
rect 11271 837 11389 871
rect 11271 803 11331 837
rect 11365 803 11389 837
rect 11271 769 11389 803
rect 11271 735 11331 769
rect 11365 735 11389 769
rect 11271 701 11389 735
rect 11271 667 11331 701
rect 11365 667 11389 701
rect 11271 633 11389 667
rect 11271 599 11331 633
rect 11365 599 11389 633
rect 11271 565 11389 599
rect 11271 531 11331 565
rect 11365 531 11389 565
rect 11271 497 11389 531
rect 7243 429 7371 463
rect 7243 395 7277 429
rect 7311 395 7371 429
rect 7243 324 7371 395
rect 11271 463 11331 497
rect 11365 463 11389 497
rect 11271 429 11389 463
rect 11271 395 11331 429
rect 11365 395 11389 429
rect 11271 324 11389 395
rect 7243 286 11389 324
rect 7243 252 7343 286
rect 7377 252 7411 286
rect 7445 252 7479 286
rect 7513 252 7547 286
rect 7581 252 7615 286
rect 7649 252 7683 286
rect 7717 252 7751 286
rect 7785 252 7819 286
rect 7853 252 7887 286
rect 7921 252 7955 286
rect 7989 252 8023 286
rect 8057 252 8091 286
rect 8125 252 8159 286
rect 8193 252 8227 286
rect 8261 252 8295 286
rect 8329 252 8363 286
rect 8397 252 8431 286
rect 8465 252 8499 286
rect 8533 252 8567 286
rect 8601 252 8635 286
rect 8669 252 8703 286
rect 8737 252 8771 286
rect 8805 252 8839 286
rect 8873 252 8907 286
rect 8941 252 8975 286
rect 9009 252 9043 286
rect 9077 252 9111 286
rect 9145 252 9179 286
rect 9213 252 9247 286
rect 9281 252 9315 286
rect 9349 252 9383 286
rect 9417 252 9451 286
rect 9485 252 9519 286
rect 9553 252 9587 286
rect 9621 252 9655 286
rect 9689 252 9723 286
rect 9757 252 9791 286
rect 9825 252 9859 286
rect 9893 252 9927 286
rect 9961 252 9995 286
rect 10029 252 10063 286
rect 10097 252 10131 286
rect 10165 252 10199 286
rect 10233 252 10267 286
rect 10301 252 10335 286
rect 10369 252 10403 286
rect 10437 252 10471 286
rect 10505 252 10539 286
rect 10573 252 10607 286
rect 10641 252 10675 286
rect 10709 252 10743 286
rect 10777 252 10811 286
rect 10845 252 10879 286
rect 10913 252 10947 286
rect 10981 252 11015 286
rect 11049 252 11083 286
rect 11117 252 11151 286
rect 11185 252 11219 286
rect 11253 252 11389 286
rect 7243 206 11389 252
<< mvpsubdiffcont >>
rect 7554 531 7792 3421
rect 8378 531 8616 3421
rect 9202 531 9440 3421
rect 10026 531 10264 3421
rect 10850 531 11088 3421
<< mvnsubdiffcont >>
rect 7353 3660 7387 3694
rect 7421 3660 7455 3694
rect 7489 3660 7523 3694
rect 7557 3660 7591 3694
rect 7625 3660 7659 3694
rect 7693 3660 7727 3694
rect 7761 3660 7795 3694
rect 7829 3660 7863 3694
rect 7897 3660 7931 3694
rect 7965 3660 7999 3694
rect 8033 3660 8067 3694
rect 8101 3660 8135 3694
rect 8169 3660 8203 3694
rect 8237 3660 8271 3694
rect 8305 3660 8339 3694
rect 8373 3660 8407 3694
rect 8441 3660 8475 3694
rect 8509 3660 8543 3694
rect 8577 3660 8611 3694
rect 8645 3660 8679 3694
rect 8713 3660 8747 3694
rect 8781 3660 8815 3694
rect 8849 3660 8883 3694
rect 8917 3660 8951 3694
rect 8985 3660 9019 3694
rect 9053 3660 9087 3694
rect 9121 3660 9155 3694
rect 9189 3660 9223 3694
rect 9257 3660 9291 3694
rect 9325 3660 9359 3694
rect 9393 3660 9427 3694
rect 9461 3660 9495 3694
rect 9529 3660 9563 3694
rect 9597 3660 9631 3694
rect 9665 3660 9699 3694
rect 9733 3660 9767 3694
rect 9801 3660 9835 3694
rect 9869 3660 9903 3694
rect 9937 3660 9971 3694
rect 10005 3660 10039 3694
rect 10073 3660 10107 3694
rect 10141 3660 10175 3694
rect 10209 3660 10243 3694
rect 10277 3660 10311 3694
rect 10345 3660 10379 3694
rect 10413 3660 10447 3694
rect 10481 3660 10515 3694
rect 10549 3660 10583 3694
rect 10617 3660 10651 3694
rect 10685 3660 10719 3694
rect 10753 3660 10787 3694
rect 10821 3660 10855 3694
rect 10889 3660 10923 3694
rect 10957 3660 10991 3694
rect 11025 3660 11059 3694
rect 11093 3660 11127 3694
rect 11161 3660 11195 3694
rect 11229 3660 11263 3694
rect 7277 3523 7311 3557
rect 7277 3455 7311 3489
rect 11331 3523 11365 3557
rect 7277 3387 7311 3421
rect 7277 3319 7311 3353
rect 7277 3251 7311 3285
rect 7277 3183 7311 3217
rect 7277 3115 7311 3149
rect 7277 3047 7311 3081
rect 7277 2979 7311 3013
rect 7277 2911 7311 2945
rect 7277 2843 7311 2877
rect 7277 2775 7311 2809
rect 7277 2707 7311 2741
rect 7277 2639 7311 2673
rect 7277 2571 7311 2605
rect 7277 2503 7311 2537
rect 7277 2435 7311 2469
rect 7277 2367 7311 2401
rect 7277 2299 7311 2333
rect 7277 2231 7311 2265
rect 7277 2163 7311 2197
rect 7277 2095 7311 2129
rect 7277 2027 7311 2061
rect 7277 1959 7311 1993
rect 7277 1891 7311 1925
rect 7277 1823 7311 1857
rect 7277 1755 7311 1789
rect 7277 1687 7311 1721
rect 7277 1619 7311 1653
rect 7277 1551 7311 1585
rect 7277 1483 7311 1517
rect 7277 1415 7311 1449
rect 7277 1347 7311 1381
rect 7277 1279 7311 1313
rect 7277 1211 7311 1245
rect 7277 1143 7311 1177
rect 7277 1075 7311 1109
rect 7277 1007 7311 1041
rect 7277 939 7311 973
rect 7277 871 7311 905
rect 7277 803 7311 837
rect 7277 735 7311 769
rect 7277 667 7311 701
rect 7277 599 7311 633
rect 7277 531 7311 565
rect 7277 463 7311 497
rect 11331 3455 11365 3489
rect 11331 3387 11365 3421
rect 11331 3319 11365 3353
rect 11331 3251 11365 3285
rect 11331 3183 11365 3217
rect 11331 3115 11365 3149
rect 11331 3047 11365 3081
rect 11331 2979 11365 3013
rect 11331 2911 11365 2945
rect 11331 2843 11365 2877
rect 11331 2775 11365 2809
rect 11331 2707 11365 2741
rect 11331 2639 11365 2673
rect 11331 2571 11365 2605
rect 11331 2503 11365 2537
rect 11331 2435 11365 2469
rect 11331 2367 11365 2401
rect 11331 2299 11365 2333
rect 11331 2231 11365 2265
rect 11331 2163 11365 2197
rect 11331 2095 11365 2129
rect 11331 2027 11365 2061
rect 11331 1959 11365 1993
rect 11331 1891 11365 1925
rect 11331 1823 11365 1857
rect 11331 1755 11365 1789
rect 11331 1687 11365 1721
rect 11331 1619 11365 1653
rect 11331 1551 11365 1585
rect 11331 1483 11365 1517
rect 11331 1415 11365 1449
rect 11331 1347 11365 1381
rect 11331 1279 11365 1313
rect 11331 1211 11365 1245
rect 11331 1143 11365 1177
rect 11331 1075 11365 1109
rect 11331 1007 11365 1041
rect 11331 939 11365 973
rect 11331 871 11365 905
rect 11331 803 11365 837
rect 11331 735 11365 769
rect 11331 667 11365 701
rect 11331 599 11365 633
rect 11331 531 11365 565
rect 7277 395 7311 429
rect 11331 463 11365 497
rect 11331 395 11365 429
rect 7343 252 7377 286
rect 7411 252 7445 286
rect 7479 252 7513 286
rect 7547 252 7581 286
rect 7615 252 7649 286
rect 7683 252 7717 286
rect 7751 252 7785 286
rect 7819 252 7853 286
rect 7887 252 7921 286
rect 7955 252 7989 286
rect 8023 252 8057 286
rect 8091 252 8125 286
rect 8159 252 8193 286
rect 8227 252 8261 286
rect 8295 252 8329 286
rect 8363 252 8397 286
rect 8431 252 8465 286
rect 8499 252 8533 286
rect 8567 252 8601 286
rect 8635 252 8669 286
rect 8703 252 8737 286
rect 8771 252 8805 286
rect 8839 252 8873 286
rect 8907 252 8941 286
rect 8975 252 9009 286
rect 9043 252 9077 286
rect 9111 252 9145 286
rect 9179 252 9213 286
rect 9247 252 9281 286
rect 9315 252 9349 286
rect 9383 252 9417 286
rect 9451 252 9485 286
rect 9519 252 9553 286
rect 9587 252 9621 286
rect 9655 252 9689 286
rect 9723 252 9757 286
rect 9791 252 9825 286
rect 9859 252 9893 286
rect 9927 252 9961 286
rect 9995 252 10029 286
rect 10063 252 10097 286
rect 10131 252 10165 286
rect 10199 252 10233 286
rect 10267 252 10301 286
rect 10335 252 10369 286
rect 10403 252 10437 286
rect 10471 252 10505 286
rect 10539 252 10573 286
rect 10607 252 10641 286
rect 10675 252 10709 286
rect 10743 252 10777 286
rect 10811 252 10845 286
rect 10879 252 10913 286
rect 10947 252 10981 286
rect 11015 252 11049 286
rect 11083 252 11117 286
rect 11151 252 11185 286
rect 11219 252 11253 286
<< mvndiode >>
rect 7935 3421 8235 3476
rect 7935 531 7966 3421
rect 8204 531 8235 3421
rect 7935 476 8235 531
rect 8759 3421 9059 3476
rect 8759 531 8790 3421
rect 9028 531 9059 3421
rect 8759 476 9059 531
rect 9583 3421 9883 3476
rect 9583 531 9614 3421
rect 9852 531 9883 3421
rect 9583 476 9883 531
rect 10407 3421 10707 3476
rect 10407 531 10438 3421
rect 10676 531 10707 3421
rect 10407 476 10707 531
<< mvndiodec >>
rect 7966 531 8204 3421
rect 8790 531 9028 3421
rect 9614 531 9852 3421
rect 10438 531 10676 3421
<< locali >>
rect 7243 3712 11389 3746
rect 7243 3678 7352 3712
rect 7386 3694 7501 3712
rect 7535 3694 7574 3712
rect 7608 3694 7646 3712
rect 7680 3694 7718 3712
rect 7752 3694 7790 3712
rect 7824 3694 7862 3712
rect 7896 3694 7934 3712
rect 7968 3694 8006 3712
rect 8040 3694 8078 3712
rect 8112 3694 8150 3712
rect 8184 3694 8222 3712
rect 8256 3694 8294 3712
rect 8328 3694 8366 3712
rect 8400 3694 8438 3712
rect 8472 3694 8510 3712
rect 8544 3694 8582 3712
rect 8616 3694 8654 3712
rect 8688 3694 8726 3712
rect 8760 3694 8798 3712
rect 8832 3694 8870 3712
rect 8904 3694 8942 3712
rect 8976 3694 9014 3712
rect 9048 3694 9086 3712
rect 9120 3694 9158 3712
rect 9192 3694 9230 3712
rect 9264 3694 9302 3712
rect 9336 3694 9374 3712
rect 9408 3694 9446 3712
rect 9480 3694 9518 3712
rect 9552 3694 9590 3712
rect 9624 3694 9662 3712
rect 9696 3694 9734 3712
rect 9768 3694 9806 3712
rect 9840 3694 9878 3712
rect 9912 3694 9950 3712
rect 9984 3694 10022 3712
rect 10056 3694 10094 3712
rect 10128 3694 10166 3712
rect 10200 3694 10238 3712
rect 10272 3694 10310 3712
rect 10344 3694 10382 3712
rect 10416 3694 10454 3712
rect 10488 3694 10526 3712
rect 10560 3694 10598 3712
rect 10632 3694 10670 3712
rect 10704 3694 10742 3712
rect 10776 3694 10814 3712
rect 10848 3694 10886 3712
rect 10920 3694 10958 3712
rect 10992 3694 11030 3712
rect 11064 3694 11102 3712
rect 11136 3694 11250 3712
rect 7243 3660 7353 3678
rect 7387 3660 7421 3694
rect 7455 3660 7489 3694
rect 7535 3678 7557 3694
rect 7608 3678 7625 3694
rect 7680 3678 7693 3694
rect 7752 3678 7761 3694
rect 7824 3678 7829 3694
rect 7896 3678 7897 3694
rect 7523 3660 7557 3678
rect 7591 3660 7625 3678
rect 7659 3660 7693 3678
rect 7727 3660 7761 3678
rect 7795 3660 7829 3678
rect 7863 3660 7897 3678
rect 7931 3678 7934 3694
rect 7999 3678 8006 3694
rect 8067 3678 8078 3694
rect 8135 3678 8150 3694
rect 8203 3678 8222 3694
rect 8271 3678 8294 3694
rect 8339 3678 8366 3694
rect 8407 3678 8438 3694
rect 7931 3660 7965 3678
rect 7999 3660 8033 3678
rect 8067 3660 8101 3678
rect 8135 3660 8169 3678
rect 8203 3660 8237 3678
rect 8271 3660 8305 3678
rect 8339 3660 8373 3678
rect 8407 3660 8441 3678
rect 8475 3660 8509 3694
rect 8544 3678 8577 3694
rect 8616 3678 8645 3694
rect 8688 3678 8713 3694
rect 8760 3678 8781 3694
rect 8832 3678 8849 3694
rect 8904 3678 8917 3694
rect 8976 3678 8985 3694
rect 9048 3678 9053 3694
rect 9120 3678 9121 3694
rect 8543 3660 8577 3678
rect 8611 3660 8645 3678
rect 8679 3660 8713 3678
rect 8747 3660 8781 3678
rect 8815 3660 8849 3678
rect 8883 3660 8917 3678
rect 8951 3660 8985 3678
rect 9019 3660 9053 3678
rect 9087 3660 9121 3678
rect 9155 3678 9158 3694
rect 9223 3678 9230 3694
rect 9291 3678 9302 3694
rect 9359 3678 9374 3694
rect 9427 3678 9446 3694
rect 9495 3678 9518 3694
rect 9563 3678 9590 3694
rect 9631 3678 9662 3694
rect 9155 3660 9189 3678
rect 9223 3660 9257 3678
rect 9291 3660 9325 3678
rect 9359 3660 9393 3678
rect 9427 3660 9461 3678
rect 9495 3660 9529 3678
rect 9563 3660 9597 3678
rect 9631 3660 9665 3678
rect 9699 3660 9733 3694
rect 9768 3678 9801 3694
rect 9840 3678 9869 3694
rect 9912 3678 9937 3694
rect 9984 3678 10005 3694
rect 10056 3678 10073 3694
rect 10128 3678 10141 3694
rect 10200 3678 10209 3694
rect 10272 3678 10277 3694
rect 10344 3678 10345 3694
rect 9767 3660 9801 3678
rect 9835 3660 9869 3678
rect 9903 3660 9937 3678
rect 9971 3660 10005 3678
rect 10039 3660 10073 3678
rect 10107 3660 10141 3678
rect 10175 3660 10209 3678
rect 10243 3660 10277 3678
rect 10311 3660 10345 3678
rect 10379 3678 10382 3694
rect 10447 3678 10454 3694
rect 10515 3678 10526 3694
rect 10583 3678 10598 3694
rect 10651 3678 10670 3694
rect 10719 3678 10742 3694
rect 10787 3678 10814 3694
rect 10855 3678 10886 3694
rect 10379 3660 10413 3678
rect 10447 3660 10481 3678
rect 10515 3660 10549 3678
rect 10583 3660 10617 3678
rect 10651 3660 10685 3678
rect 10719 3660 10753 3678
rect 10787 3660 10821 3678
rect 10855 3660 10889 3678
rect 10923 3660 10957 3694
rect 10992 3678 11025 3694
rect 11064 3678 11093 3694
rect 11136 3678 11161 3694
rect 10991 3660 11025 3678
rect 11059 3660 11093 3678
rect 11127 3660 11161 3678
rect 11195 3660 11229 3694
rect 11284 3678 11389 3712
rect 11263 3660 11389 3678
rect 7243 3628 11389 3660
rect 7243 3557 7335 3628
rect 7243 3548 7277 3557
rect 7243 3514 7274 3548
rect 7311 3523 7335 3557
rect 7308 3514 7335 3523
rect 7243 3489 7335 3514
rect 7243 3464 7277 3489
rect 7243 3430 7274 3464
rect 7311 3455 7335 3489
rect 11307 3557 11389 3628
rect 11307 3548 11331 3557
rect 11307 3514 11328 3548
rect 11365 3523 11389 3557
rect 11362 3514 11389 3523
rect 11307 3489 11389 3514
rect 7308 3430 7335 3455
rect 7243 3421 7335 3430
rect 7243 3392 7277 3421
rect 7243 3358 7274 3392
rect 7311 3387 7335 3421
rect 7308 3358 7335 3387
rect 7243 3353 7335 3358
rect 7243 3320 7277 3353
rect 7243 3286 7274 3320
rect 7311 3319 7335 3353
rect 7308 3286 7335 3319
rect 7243 3285 7335 3286
rect 7243 3251 7277 3285
rect 7311 3251 7335 3285
rect 7243 3248 7335 3251
rect 7243 3214 7274 3248
rect 7308 3217 7335 3248
rect 7243 3183 7277 3214
rect 7311 3183 7335 3217
rect 7243 3176 7335 3183
rect 7243 3142 7274 3176
rect 7308 3149 7335 3176
rect 7243 3115 7277 3142
rect 7311 3115 7335 3149
rect 7243 3104 7335 3115
rect 7243 3070 7274 3104
rect 7308 3081 7335 3104
rect 7243 3047 7277 3070
rect 7311 3047 7335 3081
rect 7243 3032 7335 3047
rect 7243 2998 7274 3032
rect 7308 3013 7335 3032
rect 7243 2979 7277 2998
rect 7311 2979 7335 3013
rect 7243 2960 7335 2979
rect 7243 2926 7274 2960
rect 7308 2945 7335 2960
rect 7243 2911 7277 2926
rect 7311 2911 7335 2945
rect 7243 2888 7335 2911
rect 7243 2854 7274 2888
rect 7308 2877 7335 2888
rect 7243 2843 7277 2854
rect 7311 2843 7335 2877
rect 7243 2816 7335 2843
rect 7243 2782 7274 2816
rect 7308 2809 7335 2816
rect 7243 2775 7277 2782
rect 7311 2775 7335 2809
rect 7243 2744 7335 2775
rect 7243 2710 7274 2744
rect 7308 2741 7335 2744
rect 7243 2707 7277 2710
rect 7311 2707 7335 2741
rect 7243 2673 7335 2707
rect 7243 2672 7277 2673
rect 7243 2638 7274 2672
rect 7311 2639 7335 2673
rect 7308 2638 7335 2639
rect 7243 2605 7335 2638
rect 7243 2600 7277 2605
rect 7243 2566 7274 2600
rect 7311 2571 7335 2605
rect 7308 2566 7335 2571
rect 7243 2537 7335 2566
rect 7243 2528 7277 2537
rect 7243 2494 7274 2528
rect 7311 2503 7335 2537
rect 7308 2494 7335 2503
rect 7243 2469 7335 2494
rect 7243 2456 7277 2469
rect 7243 2422 7274 2456
rect 7311 2435 7335 2469
rect 7308 2422 7335 2435
rect 7243 2401 7335 2422
rect 7243 2384 7277 2401
rect 7243 2350 7274 2384
rect 7311 2367 7335 2401
rect 7308 2350 7335 2367
rect 7243 2333 7335 2350
rect 7243 2312 7277 2333
rect 7243 2278 7274 2312
rect 7311 2299 7335 2333
rect 7308 2278 7335 2299
rect 7243 2265 7335 2278
rect 7243 2240 7277 2265
rect 7243 2206 7274 2240
rect 7311 2231 7335 2265
rect 7308 2206 7335 2231
rect 7243 2197 7335 2206
rect 7243 2168 7277 2197
rect 7243 2134 7274 2168
rect 7311 2163 7335 2197
rect 7308 2134 7335 2163
rect 7243 2129 7335 2134
rect 7243 2096 7277 2129
rect 7243 2062 7274 2096
rect 7311 2095 7335 2129
rect 7308 2062 7335 2095
rect 7243 2061 7335 2062
rect 7243 2027 7277 2061
rect 7311 2027 7335 2061
rect 7243 2024 7335 2027
rect 7243 1990 7274 2024
rect 7308 1993 7335 2024
rect 7243 1959 7277 1990
rect 7311 1959 7335 1993
rect 7243 1952 7335 1959
rect 7243 1918 7274 1952
rect 7308 1925 7335 1952
rect 7243 1891 7277 1918
rect 7311 1891 7335 1925
rect 7243 1880 7335 1891
rect 7243 1846 7274 1880
rect 7308 1857 7335 1880
rect 7243 1823 7277 1846
rect 7311 1823 7335 1857
rect 7243 1808 7335 1823
rect 7243 1774 7274 1808
rect 7308 1789 7335 1808
rect 7243 1755 7277 1774
rect 7311 1755 7335 1789
rect 7243 1736 7335 1755
rect 7243 1702 7274 1736
rect 7308 1721 7335 1736
rect 7243 1687 7277 1702
rect 7311 1687 7335 1721
rect 7243 1664 7335 1687
rect 7243 1630 7274 1664
rect 7308 1653 7335 1664
rect 7243 1619 7277 1630
rect 7311 1619 7335 1653
rect 7243 1592 7335 1619
rect 7243 1558 7274 1592
rect 7308 1585 7335 1592
rect 7243 1551 7277 1558
rect 7311 1551 7335 1585
rect 7243 1520 7335 1551
rect 7243 1486 7274 1520
rect 7308 1517 7335 1520
rect 7243 1483 7277 1486
rect 7311 1483 7335 1517
rect 7243 1449 7335 1483
rect 7243 1448 7277 1449
rect 7243 1414 7274 1448
rect 7311 1415 7335 1449
rect 7308 1414 7335 1415
rect 7243 1381 7335 1414
rect 7243 1376 7277 1381
rect 7243 1342 7274 1376
rect 7311 1347 7335 1381
rect 7308 1342 7335 1347
rect 7243 1313 7335 1342
rect 7243 1304 7277 1313
rect 7243 1270 7274 1304
rect 7311 1279 7335 1313
rect 7308 1270 7335 1279
rect 7243 1245 7335 1270
rect 7243 1232 7277 1245
rect 7243 1198 7274 1232
rect 7311 1211 7335 1245
rect 7308 1198 7335 1211
rect 7243 1177 7335 1198
rect 7243 1160 7277 1177
rect 7243 1126 7274 1160
rect 7311 1143 7335 1177
rect 7308 1126 7335 1143
rect 7243 1109 7335 1126
rect 7243 1088 7277 1109
rect 7243 1054 7274 1088
rect 7311 1075 7335 1109
rect 7308 1054 7335 1075
rect 7243 1041 7335 1054
rect 7243 1016 7277 1041
rect 7243 982 7274 1016
rect 7311 1007 7335 1041
rect 7308 982 7335 1007
rect 7243 973 7335 982
rect 7243 944 7277 973
rect 7243 910 7274 944
rect 7311 939 7335 973
rect 7308 910 7335 939
rect 7243 905 7335 910
rect 7243 872 7277 905
rect 7243 838 7274 872
rect 7311 871 7335 905
rect 7308 838 7335 871
rect 7243 837 7335 838
rect 7243 803 7277 837
rect 7311 803 7335 837
rect 7243 800 7335 803
rect 7243 766 7274 800
rect 7308 769 7335 800
rect 7243 735 7277 766
rect 7311 735 7335 769
rect 7243 728 7335 735
rect 7243 694 7274 728
rect 7308 701 7335 728
rect 7243 667 7277 694
rect 7311 667 7335 701
rect 7243 656 7335 667
rect 7243 622 7274 656
rect 7308 633 7335 656
rect 7243 599 7277 622
rect 7311 599 7335 633
rect 7243 565 7335 599
rect 7243 531 7277 565
rect 7311 531 7335 565
rect 7243 497 7335 531
rect 7243 463 7277 497
rect 7311 463 7335 497
rect 7523 3421 7823 3476
rect 7523 531 7554 3421
rect 7792 531 7823 3421
rect 7523 476 7823 531
rect 7935 3421 8235 3476
rect 7935 531 7966 3421
rect 8204 531 8235 3421
rect 7935 476 8235 531
rect 8347 3421 8647 3476
rect 8347 531 8378 3421
rect 8616 531 8647 3421
rect 8347 476 8647 531
rect 8759 3421 9059 3476
rect 8759 531 8790 3421
rect 9028 531 9059 3421
rect 8759 476 9059 531
rect 9171 3421 9471 3476
rect 9171 531 9202 3421
rect 9440 531 9471 3421
rect 9171 476 9471 531
rect 9583 3421 9883 3476
rect 9583 531 9614 3421
rect 9852 531 9883 3421
rect 9583 476 9883 531
rect 9995 3421 10295 3476
rect 9995 531 10026 3421
rect 10264 531 10295 3421
rect 9995 476 10295 531
rect 10407 3421 10707 3476
rect 10407 531 10438 3421
rect 10676 531 10707 3421
rect 10407 476 10707 531
rect 10819 3421 11119 3476
rect 10819 531 10850 3421
rect 11088 531 11119 3421
rect 10819 476 11119 531
rect 11307 3464 11331 3489
rect 11307 3430 11328 3464
rect 11365 3455 11389 3489
rect 11362 3430 11389 3455
rect 11307 3421 11389 3430
rect 11307 3392 11331 3421
rect 11307 3358 11328 3392
rect 11365 3387 11389 3421
rect 11362 3358 11389 3387
rect 11307 3353 11389 3358
rect 11307 3320 11331 3353
rect 11307 3286 11328 3320
rect 11365 3319 11389 3353
rect 11362 3286 11389 3319
rect 11307 3285 11389 3286
rect 11307 3251 11331 3285
rect 11365 3251 11389 3285
rect 11307 3248 11389 3251
rect 11307 3214 11328 3248
rect 11362 3217 11389 3248
rect 11307 3183 11331 3214
rect 11365 3183 11389 3217
rect 11307 3176 11389 3183
rect 11307 3142 11328 3176
rect 11362 3149 11389 3176
rect 11307 3115 11331 3142
rect 11365 3115 11389 3149
rect 11307 3104 11389 3115
rect 11307 3070 11328 3104
rect 11362 3081 11389 3104
rect 11307 3047 11331 3070
rect 11365 3047 11389 3081
rect 11307 3032 11389 3047
rect 11307 2998 11328 3032
rect 11362 3013 11389 3032
rect 11307 2979 11331 2998
rect 11365 2979 11389 3013
rect 11307 2960 11389 2979
rect 11307 2926 11328 2960
rect 11362 2945 11389 2960
rect 11307 2911 11331 2926
rect 11365 2911 11389 2945
rect 11307 2888 11389 2911
rect 11307 2854 11328 2888
rect 11362 2877 11389 2888
rect 11307 2843 11331 2854
rect 11365 2843 11389 2877
rect 11307 2816 11389 2843
rect 11307 2782 11328 2816
rect 11362 2809 11389 2816
rect 11307 2775 11331 2782
rect 11365 2775 11389 2809
rect 11307 2744 11389 2775
rect 11307 2710 11328 2744
rect 11362 2741 11389 2744
rect 11307 2707 11331 2710
rect 11365 2707 11389 2741
rect 11307 2673 11389 2707
rect 11307 2672 11331 2673
rect 11307 2638 11328 2672
rect 11365 2639 11389 2673
rect 11362 2638 11389 2639
rect 11307 2605 11389 2638
rect 11307 2600 11331 2605
rect 11307 2566 11328 2600
rect 11365 2571 11389 2605
rect 11362 2566 11389 2571
rect 11307 2537 11389 2566
rect 11307 2528 11331 2537
rect 11307 2494 11328 2528
rect 11365 2503 11389 2537
rect 11362 2494 11389 2503
rect 11307 2469 11389 2494
rect 11307 2456 11331 2469
rect 11307 2422 11328 2456
rect 11365 2435 11389 2469
rect 11362 2422 11389 2435
rect 11307 2401 11389 2422
rect 11307 2384 11331 2401
rect 11307 2350 11328 2384
rect 11365 2367 11389 2401
rect 11362 2350 11389 2367
rect 11307 2333 11389 2350
rect 11307 2312 11331 2333
rect 11307 2278 11328 2312
rect 11365 2299 11389 2333
rect 11362 2278 11389 2299
rect 11307 2265 11389 2278
rect 11307 2240 11331 2265
rect 11307 2206 11328 2240
rect 11365 2231 11389 2265
rect 11362 2206 11389 2231
rect 11307 2197 11389 2206
rect 11307 2168 11331 2197
rect 11307 2134 11328 2168
rect 11365 2163 11389 2197
rect 11362 2134 11389 2163
rect 11307 2129 11389 2134
rect 11307 2096 11331 2129
rect 11307 2062 11328 2096
rect 11365 2095 11389 2129
rect 11362 2062 11389 2095
rect 11307 2061 11389 2062
rect 11307 2027 11331 2061
rect 11365 2027 11389 2061
rect 11307 2024 11389 2027
rect 11307 1990 11328 2024
rect 11362 1993 11389 2024
rect 11307 1959 11331 1990
rect 11365 1959 11389 1993
rect 11307 1952 11389 1959
rect 11307 1918 11328 1952
rect 11362 1925 11389 1952
rect 11307 1891 11331 1918
rect 11365 1891 11389 1925
rect 11307 1880 11389 1891
rect 11307 1846 11328 1880
rect 11362 1857 11389 1880
rect 11307 1823 11331 1846
rect 11365 1823 11389 1857
rect 11307 1808 11389 1823
rect 11307 1774 11328 1808
rect 11362 1789 11389 1808
rect 11307 1755 11331 1774
rect 11365 1755 11389 1789
rect 11307 1736 11389 1755
rect 11307 1702 11328 1736
rect 11362 1721 11389 1736
rect 11307 1687 11331 1702
rect 11365 1687 11389 1721
rect 11307 1664 11389 1687
rect 11307 1630 11328 1664
rect 11362 1653 11389 1664
rect 11307 1619 11331 1630
rect 11365 1619 11389 1653
rect 11307 1592 11389 1619
rect 11307 1558 11328 1592
rect 11362 1585 11389 1592
rect 11307 1551 11331 1558
rect 11365 1551 11389 1585
rect 11307 1520 11389 1551
rect 11307 1486 11328 1520
rect 11362 1517 11389 1520
rect 11307 1483 11331 1486
rect 11365 1483 11389 1517
rect 11307 1449 11389 1483
rect 11307 1448 11331 1449
rect 11307 1414 11328 1448
rect 11365 1415 11389 1449
rect 11362 1414 11389 1415
rect 11307 1381 11389 1414
rect 11307 1376 11331 1381
rect 11307 1342 11328 1376
rect 11365 1347 11389 1381
rect 11362 1342 11389 1347
rect 11307 1313 11389 1342
rect 11307 1304 11331 1313
rect 11307 1270 11328 1304
rect 11365 1279 11389 1313
rect 11362 1270 11389 1279
rect 11307 1245 11389 1270
rect 11307 1232 11331 1245
rect 11307 1198 11328 1232
rect 11365 1211 11389 1245
rect 11362 1198 11389 1211
rect 11307 1177 11389 1198
rect 11307 1160 11331 1177
rect 11307 1126 11328 1160
rect 11365 1143 11389 1177
rect 11362 1126 11389 1143
rect 11307 1109 11389 1126
rect 11307 1088 11331 1109
rect 11307 1054 11328 1088
rect 11365 1075 11389 1109
rect 11362 1054 11389 1075
rect 11307 1041 11389 1054
rect 11307 1016 11331 1041
rect 11307 982 11328 1016
rect 11365 1007 11389 1041
rect 11362 982 11389 1007
rect 11307 973 11389 982
rect 11307 944 11331 973
rect 11307 910 11328 944
rect 11365 939 11389 973
rect 11362 910 11389 939
rect 11307 905 11389 910
rect 11307 872 11331 905
rect 11307 838 11328 872
rect 11365 871 11389 905
rect 11362 838 11389 871
rect 11307 837 11389 838
rect 11307 803 11331 837
rect 11365 803 11389 837
rect 11307 800 11389 803
rect 11307 766 11328 800
rect 11362 769 11389 800
rect 11307 735 11331 766
rect 11365 735 11389 769
rect 11307 728 11389 735
rect 11307 694 11328 728
rect 11362 701 11389 728
rect 11307 667 11331 694
rect 11365 667 11389 701
rect 11307 656 11389 667
rect 11307 622 11328 656
rect 11362 633 11389 656
rect 11307 599 11331 622
rect 11365 599 11389 633
rect 11307 565 11389 599
rect 11307 531 11331 565
rect 11365 531 11389 565
rect 11307 497 11389 531
rect 7243 429 7335 463
rect 7243 395 7277 429
rect 7311 395 7335 429
rect 7243 316 7335 395
rect 11307 463 11331 497
rect 11365 463 11389 497
rect 11307 429 11389 463
rect 11307 395 11331 429
rect 11365 395 11389 429
rect 11307 316 11389 395
rect 7243 286 11389 316
rect 7243 252 7343 286
rect 7377 252 7411 286
rect 7445 252 7479 286
rect 7513 252 7547 286
rect 7581 252 7615 286
rect 7649 252 7683 286
rect 7717 252 7751 286
rect 7785 252 7819 286
rect 7853 252 7887 286
rect 7921 252 7955 286
rect 7989 252 8023 286
rect 8057 252 8091 286
rect 8125 252 8159 286
rect 8193 252 8227 286
rect 8261 252 8295 286
rect 8329 252 8363 286
rect 8397 252 8431 286
rect 8465 252 8499 286
rect 8533 252 8567 286
rect 8601 252 8635 286
rect 8669 252 8703 286
rect 8737 252 8771 286
rect 8805 252 8839 286
rect 8873 252 8907 286
rect 8941 252 8975 286
rect 9009 252 9043 286
rect 9077 252 9111 286
rect 9145 252 9179 286
rect 9213 252 9247 286
rect 9281 252 9315 286
rect 9349 252 9383 286
rect 9417 252 9451 286
rect 9485 252 9519 286
rect 9553 252 9587 286
rect 9621 252 9655 286
rect 9689 252 9723 286
rect 9757 252 9791 286
rect 9825 252 9859 286
rect 9893 252 9927 286
rect 9961 252 9995 286
rect 10029 252 10063 286
rect 10097 252 10131 286
rect 10165 252 10199 286
rect 10233 252 10267 286
rect 10301 252 10335 286
rect 10369 252 10403 286
rect 10437 252 10471 286
rect 10505 252 10539 286
rect 10573 252 10607 286
rect 10641 252 10675 286
rect 10709 252 10743 286
rect 10777 252 10811 286
rect 10845 252 10879 286
rect 10913 252 10947 286
rect 10981 252 11015 286
rect 11049 252 11083 286
rect 11117 252 11151 286
rect 11185 252 11219 286
rect 11253 252 11389 286
rect 7243 206 11389 252
<< viali >>
rect 7352 3694 7386 3712
rect 7501 3694 7535 3712
rect 7574 3694 7608 3712
rect 7646 3694 7680 3712
rect 7718 3694 7752 3712
rect 7790 3694 7824 3712
rect 7862 3694 7896 3712
rect 7934 3694 7968 3712
rect 8006 3694 8040 3712
rect 8078 3694 8112 3712
rect 8150 3694 8184 3712
rect 8222 3694 8256 3712
rect 8294 3694 8328 3712
rect 8366 3694 8400 3712
rect 8438 3694 8472 3712
rect 8510 3694 8544 3712
rect 8582 3694 8616 3712
rect 8654 3694 8688 3712
rect 8726 3694 8760 3712
rect 8798 3694 8832 3712
rect 8870 3694 8904 3712
rect 8942 3694 8976 3712
rect 9014 3694 9048 3712
rect 9086 3694 9120 3712
rect 9158 3694 9192 3712
rect 9230 3694 9264 3712
rect 9302 3694 9336 3712
rect 9374 3694 9408 3712
rect 9446 3694 9480 3712
rect 9518 3694 9552 3712
rect 9590 3694 9624 3712
rect 9662 3694 9696 3712
rect 9734 3694 9768 3712
rect 9806 3694 9840 3712
rect 9878 3694 9912 3712
rect 9950 3694 9984 3712
rect 10022 3694 10056 3712
rect 10094 3694 10128 3712
rect 10166 3694 10200 3712
rect 10238 3694 10272 3712
rect 10310 3694 10344 3712
rect 10382 3694 10416 3712
rect 10454 3694 10488 3712
rect 10526 3694 10560 3712
rect 10598 3694 10632 3712
rect 10670 3694 10704 3712
rect 10742 3694 10776 3712
rect 10814 3694 10848 3712
rect 10886 3694 10920 3712
rect 10958 3694 10992 3712
rect 11030 3694 11064 3712
rect 11102 3694 11136 3712
rect 11250 3694 11284 3712
rect 7352 3678 7353 3694
rect 7353 3678 7386 3694
rect 7501 3678 7523 3694
rect 7523 3678 7535 3694
rect 7574 3678 7591 3694
rect 7591 3678 7608 3694
rect 7646 3678 7659 3694
rect 7659 3678 7680 3694
rect 7718 3678 7727 3694
rect 7727 3678 7752 3694
rect 7790 3678 7795 3694
rect 7795 3678 7824 3694
rect 7862 3678 7863 3694
rect 7863 3678 7896 3694
rect 7934 3678 7965 3694
rect 7965 3678 7968 3694
rect 8006 3678 8033 3694
rect 8033 3678 8040 3694
rect 8078 3678 8101 3694
rect 8101 3678 8112 3694
rect 8150 3678 8169 3694
rect 8169 3678 8184 3694
rect 8222 3678 8237 3694
rect 8237 3678 8256 3694
rect 8294 3678 8305 3694
rect 8305 3678 8328 3694
rect 8366 3678 8373 3694
rect 8373 3678 8400 3694
rect 8438 3678 8441 3694
rect 8441 3678 8472 3694
rect 8510 3678 8543 3694
rect 8543 3678 8544 3694
rect 8582 3678 8611 3694
rect 8611 3678 8616 3694
rect 8654 3678 8679 3694
rect 8679 3678 8688 3694
rect 8726 3678 8747 3694
rect 8747 3678 8760 3694
rect 8798 3678 8815 3694
rect 8815 3678 8832 3694
rect 8870 3678 8883 3694
rect 8883 3678 8904 3694
rect 8942 3678 8951 3694
rect 8951 3678 8976 3694
rect 9014 3678 9019 3694
rect 9019 3678 9048 3694
rect 9086 3678 9087 3694
rect 9087 3678 9120 3694
rect 9158 3678 9189 3694
rect 9189 3678 9192 3694
rect 9230 3678 9257 3694
rect 9257 3678 9264 3694
rect 9302 3678 9325 3694
rect 9325 3678 9336 3694
rect 9374 3678 9393 3694
rect 9393 3678 9408 3694
rect 9446 3678 9461 3694
rect 9461 3678 9480 3694
rect 9518 3678 9529 3694
rect 9529 3678 9552 3694
rect 9590 3678 9597 3694
rect 9597 3678 9624 3694
rect 9662 3678 9665 3694
rect 9665 3678 9696 3694
rect 9734 3678 9767 3694
rect 9767 3678 9768 3694
rect 9806 3678 9835 3694
rect 9835 3678 9840 3694
rect 9878 3678 9903 3694
rect 9903 3678 9912 3694
rect 9950 3678 9971 3694
rect 9971 3678 9984 3694
rect 10022 3678 10039 3694
rect 10039 3678 10056 3694
rect 10094 3678 10107 3694
rect 10107 3678 10128 3694
rect 10166 3678 10175 3694
rect 10175 3678 10200 3694
rect 10238 3678 10243 3694
rect 10243 3678 10272 3694
rect 10310 3678 10311 3694
rect 10311 3678 10344 3694
rect 10382 3678 10413 3694
rect 10413 3678 10416 3694
rect 10454 3678 10481 3694
rect 10481 3678 10488 3694
rect 10526 3678 10549 3694
rect 10549 3678 10560 3694
rect 10598 3678 10617 3694
rect 10617 3678 10632 3694
rect 10670 3678 10685 3694
rect 10685 3678 10704 3694
rect 10742 3678 10753 3694
rect 10753 3678 10776 3694
rect 10814 3678 10821 3694
rect 10821 3678 10848 3694
rect 10886 3678 10889 3694
rect 10889 3678 10920 3694
rect 10958 3678 10991 3694
rect 10991 3678 10992 3694
rect 11030 3678 11059 3694
rect 11059 3678 11064 3694
rect 11102 3678 11127 3694
rect 11127 3678 11136 3694
rect 11250 3678 11263 3694
rect 11263 3678 11284 3694
rect 7274 3523 7277 3548
rect 7277 3523 7308 3548
rect 7274 3514 7308 3523
rect 7274 3455 7277 3464
rect 7277 3455 7308 3464
rect 11328 3523 11331 3548
rect 11331 3523 11362 3548
rect 11328 3514 11362 3523
rect 7274 3430 7308 3455
rect 7274 3387 7277 3392
rect 7277 3387 7308 3392
rect 7274 3358 7308 3387
rect 7274 3319 7277 3320
rect 7277 3319 7308 3320
rect 7274 3286 7308 3319
rect 7274 3217 7308 3248
rect 7274 3214 7277 3217
rect 7277 3214 7308 3217
rect 7274 3149 7308 3176
rect 7274 3142 7277 3149
rect 7277 3142 7308 3149
rect 7274 3081 7308 3104
rect 7274 3070 7277 3081
rect 7277 3070 7308 3081
rect 7274 3013 7308 3032
rect 7274 2998 7277 3013
rect 7277 2998 7308 3013
rect 7274 2945 7308 2960
rect 7274 2926 7277 2945
rect 7277 2926 7308 2945
rect 7274 2877 7308 2888
rect 7274 2854 7277 2877
rect 7277 2854 7308 2877
rect 7274 2809 7308 2816
rect 7274 2782 7277 2809
rect 7277 2782 7308 2809
rect 7274 2741 7308 2744
rect 7274 2710 7277 2741
rect 7277 2710 7308 2741
rect 7274 2639 7277 2672
rect 7277 2639 7308 2672
rect 7274 2638 7308 2639
rect 7274 2571 7277 2600
rect 7277 2571 7308 2600
rect 7274 2566 7308 2571
rect 7274 2503 7277 2528
rect 7277 2503 7308 2528
rect 7274 2494 7308 2503
rect 7274 2435 7277 2456
rect 7277 2435 7308 2456
rect 7274 2422 7308 2435
rect 7274 2367 7277 2384
rect 7277 2367 7308 2384
rect 7274 2350 7308 2367
rect 7274 2299 7277 2312
rect 7277 2299 7308 2312
rect 7274 2278 7308 2299
rect 7274 2231 7277 2240
rect 7277 2231 7308 2240
rect 7274 2206 7308 2231
rect 7274 2163 7277 2168
rect 7277 2163 7308 2168
rect 7274 2134 7308 2163
rect 7274 2095 7277 2096
rect 7277 2095 7308 2096
rect 7274 2062 7308 2095
rect 7274 1993 7308 2024
rect 7274 1990 7277 1993
rect 7277 1990 7308 1993
rect 7274 1925 7308 1952
rect 7274 1918 7277 1925
rect 7277 1918 7308 1925
rect 7274 1857 7308 1880
rect 7274 1846 7277 1857
rect 7277 1846 7308 1857
rect 7274 1789 7308 1808
rect 7274 1774 7277 1789
rect 7277 1774 7308 1789
rect 7274 1721 7308 1736
rect 7274 1702 7277 1721
rect 7277 1702 7308 1721
rect 7274 1653 7308 1664
rect 7274 1630 7277 1653
rect 7277 1630 7308 1653
rect 7274 1585 7308 1592
rect 7274 1558 7277 1585
rect 7277 1558 7308 1585
rect 7274 1517 7308 1520
rect 7274 1486 7277 1517
rect 7277 1486 7308 1517
rect 7274 1415 7277 1448
rect 7277 1415 7308 1448
rect 7274 1414 7308 1415
rect 7274 1347 7277 1376
rect 7277 1347 7308 1376
rect 7274 1342 7308 1347
rect 7274 1279 7277 1304
rect 7277 1279 7308 1304
rect 7274 1270 7308 1279
rect 7274 1211 7277 1232
rect 7277 1211 7308 1232
rect 7274 1198 7308 1211
rect 7274 1143 7277 1160
rect 7277 1143 7308 1160
rect 7274 1126 7308 1143
rect 7274 1075 7277 1088
rect 7277 1075 7308 1088
rect 7274 1054 7308 1075
rect 7274 1007 7277 1016
rect 7277 1007 7308 1016
rect 7274 982 7308 1007
rect 7274 939 7277 944
rect 7277 939 7308 944
rect 7274 910 7308 939
rect 7274 871 7277 872
rect 7277 871 7308 872
rect 7274 838 7308 871
rect 7274 769 7308 800
rect 7274 766 7277 769
rect 7277 766 7308 769
rect 7274 701 7308 728
rect 7274 694 7277 701
rect 7277 694 7308 701
rect 7274 633 7308 656
rect 7274 622 7277 633
rect 7277 622 7308 633
rect 7584 3303 7618 3337
rect 7656 3303 7690 3337
rect 7728 3303 7762 3337
rect 7584 3207 7618 3241
rect 7656 3207 7690 3241
rect 7728 3207 7762 3241
rect 7584 3111 7618 3145
rect 7656 3111 7690 3145
rect 7728 3111 7762 3145
rect 7584 3015 7618 3049
rect 7656 3015 7690 3049
rect 7728 3015 7762 3049
rect 7584 2919 7618 2953
rect 7656 2919 7690 2953
rect 7728 2919 7762 2953
rect 7584 2823 7618 2857
rect 7656 2823 7690 2857
rect 7728 2823 7762 2857
rect 7584 2727 7618 2761
rect 7656 2727 7690 2761
rect 7728 2727 7762 2761
rect 7584 2631 7618 2665
rect 7656 2631 7690 2665
rect 7728 2631 7762 2665
rect 7584 2535 7618 2569
rect 7656 2535 7690 2569
rect 7728 2535 7762 2569
rect 7584 2439 7618 2473
rect 7656 2439 7690 2473
rect 7728 2439 7762 2473
rect 7584 2343 7618 2377
rect 7656 2343 7690 2377
rect 7728 2343 7762 2377
rect 7584 2247 7618 2281
rect 7656 2247 7690 2281
rect 7728 2247 7762 2281
rect 7584 2151 7618 2185
rect 7656 2151 7690 2185
rect 7728 2151 7762 2185
rect 7584 2055 7618 2089
rect 7656 2055 7690 2089
rect 7728 2055 7762 2089
rect 7584 1959 7618 1993
rect 7656 1959 7690 1993
rect 7728 1959 7762 1993
rect 7584 1863 7618 1897
rect 7656 1863 7690 1897
rect 7728 1863 7762 1897
rect 7584 1767 7618 1801
rect 7656 1767 7690 1801
rect 7728 1767 7762 1801
rect 7584 1671 7618 1705
rect 7656 1671 7690 1705
rect 7728 1671 7762 1705
rect 7584 1575 7618 1609
rect 7656 1575 7690 1609
rect 7728 1575 7762 1609
rect 7584 1479 7618 1513
rect 7656 1479 7690 1513
rect 7728 1479 7762 1513
rect 7584 1383 7618 1417
rect 7656 1383 7690 1417
rect 7728 1383 7762 1417
rect 7584 1287 7618 1321
rect 7656 1287 7690 1321
rect 7728 1287 7762 1321
rect 7584 1191 7618 1225
rect 7656 1191 7690 1225
rect 7728 1191 7762 1225
rect 7584 1095 7618 1129
rect 7656 1095 7690 1129
rect 7728 1095 7762 1129
rect 7584 999 7618 1033
rect 7656 999 7690 1033
rect 7728 999 7762 1033
rect 7584 903 7618 937
rect 7656 903 7690 937
rect 7728 903 7762 937
rect 7584 807 7618 841
rect 7656 807 7690 841
rect 7728 807 7762 841
rect 7584 711 7618 745
rect 7656 711 7690 745
rect 7728 711 7762 745
rect 7584 615 7618 649
rect 7656 615 7690 649
rect 7728 615 7762 649
rect 7996 3303 8030 3337
rect 8068 3303 8102 3337
rect 8140 3303 8174 3337
rect 7996 3207 8030 3241
rect 8068 3207 8102 3241
rect 8140 3207 8174 3241
rect 7996 3111 8030 3145
rect 8068 3111 8102 3145
rect 8140 3111 8174 3145
rect 7996 3015 8030 3049
rect 8068 3015 8102 3049
rect 8140 3015 8174 3049
rect 7996 2919 8030 2953
rect 8068 2919 8102 2953
rect 8140 2919 8174 2953
rect 7996 2823 8030 2857
rect 8068 2823 8102 2857
rect 8140 2823 8174 2857
rect 7996 2727 8030 2761
rect 8068 2727 8102 2761
rect 8140 2727 8174 2761
rect 7996 2631 8030 2665
rect 8068 2631 8102 2665
rect 8140 2631 8174 2665
rect 7996 2535 8030 2569
rect 8068 2535 8102 2569
rect 8140 2535 8174 2569
rect 7996 2439 8030 2473
rect 8068 2439 8102 2473
rect 8140 2439 8174 2473
rect 7996 2343 8030 2377
rect 8068 2343 8102 2377
rect 8140 2343 8174 2377
rect 7996 2247 8030 2281
rect 8068 2247 8102 2281
rect 8140 2247 8174 2281
rect 7996 2151 8030 2185
rect 8068 2151 8102 2185
rect 8140 2151 8174 2185
rect 7996 2055 8030 2089
rect 8068 2055 8102 2089
rect 8140 2055 8174 2089
rect 7996 1959 8030 1993
rect 8068 1959 8102 1993
rect 8140 1959 8174 1993
rect 7996 1863 8030 1897
rect 8068 1863 8102 1897
rect 8140 1863 8174 1897
rect 7996 1767 8030 1801
rect 8068 1767 8102 1801
rect 8140 1767 8174 1801
rect 7996 1671 8030 1705
rect 8068 1671 8102 1705
rect 8140 1671 8174 1705
rect 7996 1575 8030 1609
rect 8068 1575 8102 1609
rect 8140 1575 8174 1609
rect 7996 1479 8030 1513
rect 8068 1479 8102 1513
rect 8140 1479 8174 1513
rect 7996 1383 8030 1417
rect 8068 1383 8102 1417
rect 8140 1383 8174 1417
rect 7996 1287 8030 1321
rect 8068 1287 8102 1321
rect 8140 1287 8174 1321
rect 7996 1191 8030 1225
rect 8068 1191 8102 1225
rect 8140 1191 8174 1225
rect 7996 1095 8030 1129
rect 8068 1095 8102 1129
rect 8140 1095 8174 1129
rect 7996 999 8030 1033
rect 8068 999 8102 1033
rect 8140 999 8174 1033
rect 7996 903 8030 937
rect 8068 903 8102 937
rect 8140 903 8174 937
rect 7996 807 8030 841
rect 8068 807 8102 841
rect 8140 807 8174 841
rect 7996 711 8030 745
rect 8068 711 8102 745
rect 8140 711 8174 745
rect 7996 615 8030 649
rect 8068 615 8102 649
rect 8140 615 8174 649
rect 8408 3303 8442 3337
rect 8480 3303 8514 3337
rect 8552 3303 8586 3337
rect 8408 3207 8442 3241
rect 8480 3207 8514 3241
rect 8552 3207 8586 3241
rect 8408 3111 8442 3145
rect 8480 3111 8514 3145
rect 8552 3111 8586 3145
rect 8408 3015 8442 3049
rect 8480 3015 8514 3049
rect 8552 3015 8586 3049
rect 8408 2919 8442 2953
rect 8480 2919 8514 2953
rect 8552 2919 8586 2953
rect 8408 2823 8442 2857
rect 8480 2823 8514 2857
rect 8552 2823 8586 2857
rect 8408 2727 8442 2761
rect 8480 2727 8514 2761
rect 8552 2727 8586 2761
rect 8408 2631 8442 2665
rect 8480 2631 8514 2665
rect 8552 2631 8586 2665
rect 8408 2535 8442 2569
rect 8480 2535 8514 2569
rect 8552 2535 8586 2569
rect 8408 2439 8442 2473
rect 8480 2439 8514 2473
rect 8552 2439 8586 2473
rect 8408 2343 8442 2377
rect 8480 2343 8514 2377
rect 8552 2343 8586 2377
rect 8408 2247 8442 2281
rect 8480 2247 8514 2281
rect 8552 2247 8586 2281
rect 8408 2151 8442 2185
rect 8480 2151 8514 2185
rect 8552 2151 8586 2185
rect 8408 2055 8442 2089
rect 8480 2055 8514 2089
rect 8552 2055 8586 2089
rect 8408 1959 8442 1993
rect 8480 1959 8514 1993
rect 8552 1959 8586 1993
rect 8408 1863 8442 1897
rect 8480 1863 8514 1897
rect 8552 1863 8586 1897
rect 8408 1767 8442 1801
rect 8480 1767 8514 1801
rect 8552 1767 8586 1801
rect 8408 1671 8442 1705
rect 8480 1671 8514 1705
rect 8552 1671 8586 1705
rect 8408 1575 8442 1609
rect 8480 1575 8514 1609
rect 8552 1575 8586 1609
rect 8408 1479 8442 1513
rect 8480 1479 8514 1513
rect 8552 1479 8586 1513
rect 8408 1383 8442 1417
rect 8480 1383 8514 1417
rect 8552 1383 8586 1417
rect 8408 1287 8442 1321
rect 8480 1287 8514 1321
rect 8552 1287 8586 1321
rect 8408 1191 8442 1225
rect 8480 1191 8514 1225
rect 8552 1191 8586 1225
rect 8408 1095 8442 1129
rect 8480 1095 8514 1129
rect 8552 1095 8586 1129
rect 8408 999 8442 1033
rect 8480 999 8514 1033
rect 8552 999 8586 1033
rect 8408 903 8442 937
rect 8480 903 8514 937
rect 8552 903 8586 937
rect 8408 807 8442 841
rect 8480 807 8514 841
rect 8552 807 8586 841
rect 8408 711 8442 745
rect 8480 711 8514 745
rect 8552 711 8586 745
rect 8408 615 8442 649
rect 8480 615 8514 649
rect 8552 615 8586 649
rect 8820 3303 8854 3337
rect 8892 3303 8926 3337
rect 8964 3303 8998 3337
rect 8820 3207 8854 3241
rect 8892 3207 8926 3241
rect 8964 3207 8998 3241
rect 8820 3111 8854 3145
rect 8892 3111 8926 3145
rect 8964 3111 8998 3145
rect 8820 3015 8854 3049
rect 8892 3015 8926 3049
rect 8964 3015 8998 3049
rect 8820 2919 8854 2953
rect 8892 2919 8926 2953
rect 8964 2919 8998 2953
rect 8820 2823 8854 2857
rect 8892 2823 8926 2857
rect 8964 2823 8998 2857
rect 8820 2727 8854 2761
rect 8892 2727 8926 2761
rect 8964 2727 8998 2761
rect 8820 2631 8854 2665
rect 8892 2631 8926 2665
rect 8964 2631 8998 2665
rect 8820 2535 8854 2569
rect 8892 2535 8926 2569
rect 8964 2535 8998 2569
rect 8820 2439 8854 2473
rect 8892 2439 8926 2473
rect 8964 2439 8998 2473
rect 8820 2343 8854 2377
rect 8892 2343 8926 2377
rect 8964 2343 8998 2377
rect 8820 2247 8854 2281
rect 8892 2247 8926 2281
rect 8964 2247 8998 2281
rect 8820 2151 8854 2185
rect 8892 2151 8926 2185
rect 8964 2151 8998 2185
rect 8820 2055 8854 2089
rect 8892 2055 8926 2089
rect 8964 2055 8998 2089
rect 8820 1959 8854 1993
rect 8892 1959 8926 1993
rect 8964 1959 8998 1993
rect 8820 1863 8854 1897
rect 8892 1863 8926 1897
rect 8964 1863 8998 1897
rect 8820 1767 8854 1801
rect 8892 1767 8926 1801
rect 8964 1767 8998 1801
rect 8820 1671 8854 1705
rect 8892 1671 8926 1705
rect 8964 1671 8998 1705
rect 8820 1575 8854 1609
rect 8892 1575 8926 1609
rect 8964 1575 8998 1609
rect 8820 1479 8854 1513
rect 8892 1479 8926 1513
rect 8964 1479 8998 1513
rect 8820 1383 8854 1417
rect 8892 1383 8926 1417
rect 8964 1383 8998 1417
rect 8820 1287 8854 1321
rect 8892 1287 8926 1321
rect 8964 1287 8998 1321
rect 8820 1191 8854 1225
rect 8892 1191 8926 1225
rect 8964 1191 8998 1225
rect 8820 1095 8854 1129
rect 8892 1095 8926 1129
rect 8964 1095 8998 1129
rect 8820 999 8854 1033
rect 8892 999 8926 1033
rect 8964 999 8998 1033
rect 8820 903 8854 937
rect 8892 903 8926 937
rect 8964 903 8998 937
rect 8820 807 8854 841
rect 8892 807 8926 841
rect 8964 807 8998 841
rect 8820 711 8854 745
rect 8892 711 8926 745
rect 8964 711 8998 745
rect 8820 615 8854 649
rect 8892 615 8926 649
rect 8964 615 8998 649
rect 9232 3303 9266 3337
rect 9304 3303 9338 3337
rect 9376 3303 9410 3337
rect 9232 3207 9266 3241
rect 9304 3207 9338 3241
rect 9376 3207 9410 3241
rect 9232 3111 9266 3145
rect 9304 3111 9338 3145
rect 9376 3111 9410 3145
rect 9232 3015 9266 3049
rect 9304 3015 9338 3049
rect 9376 3015 9410 3049
rect 9232 2919 9266 2953
rect 9304 2919 9338 2953
rect 9376 2919 9410 2953
rect 9232 2823 9266 2857
rect 9304 2823 9338 2857
rect 9376 2823 9410 2857
rect 9232 2727 9266 2761
rect 9304 2727 9338 2761
rect 9376 2727 9410 2761
rect 9232 2631 9266 2665
rect 9304 2631 9338 2665
rect 9376 2631 9410 2665
rect 9232 2535 9266 2569
rect 9304 2535 9338 2569
rect 9376 2535 9410 2569
rect 9232 2439 9266 2473
rect 9304 2439 9338 2473
rect 9376 2439 9410 2473
rect 9232 2343 9266 2377
rect 9304 2343 9338 2377
rect 9376 2343 9410 2377
rect 9232 2247 9266 2281
rect 9304 2247 9338 2281
rect 9376 2247 9410 2281
rect 9232 2151 9266 2185
rect 9304 2151 9338 2185
rect 9376 2151 9410 2185
rect 9232 2055 9266 2089
rect 9304 2055 9338 2089
rect 9376 2055 9410 2089
rect 9232 1959 9266 1993
rect 9304 1959 9338 1993
rect 9376 1959 9410 1993
rect 9232 1863 9266 1897
rect 9304 1863 9338 1897
rect 9376 1863 9410 1897
rect 9232 1767 9266 1801
rect 9304 1767 9338 1801
rect 9376 1767 9410 1801
rect 9232 1671 9266 1705
rect 9304 1671 9338 1705
rect 9376 1671 9410 1705
rect 9232 1575 9266 1609
rect 9304 1575 9338 1609
rect 9376 1575 9410 1609
rect 9232 1479 9266 1513
rect 9304 1479 9338 1513
rect 9376 1479 9410 1513
rect 9232 1383 9266 1417
rect 9304 1383 9338 1417
rect 9376 1383 9410 1417
rect 9232 1287 9266 1321
rect 9304 1287 9338 1321
rect 9376 1287 9410 1321
rect 9232 1191 9266 1225
rect 9304 1191 9338 1225
rect 9376 1191 9410 1225
rect 9232 1095 9266 1129
rect 9304 1095 9338 1129
rect 9376 1095 9410 1129
rect 9232 999 9266 1033
rect 9304 999 9338 1033
rect 9376 999 9410 1033
rect 9232 903 9266 937
rect 9304 903 9338 937
rect 9376 903 9410 937
rect 9232 807 9266 841
rect 9304 807 9338 841
rect 9376 807 9410 841
rect 9232 711 9266 745
rect 9304 711 9338 745
rect 9376 711 9410 745
rect 9232 615 9266 649
rect 9304 615 9338 649
rect 9376 615 9410 649
rect 9644 3303 9678 3337
rect 9716 3303 9750 3337
rect 9788 3303 9822 3337
rect 9644 3207 9678 3241
rect 9716 3207 9750 3241
rect 9788 3207 9822 3241
rect 9644 3111 9678 3145
rect 9716 3111 9750 3145
rect 9788 3111 9822 3145
rect 9644 3015 9678 3049
rect 9716 3015 9750 3049
rect 9788 3015 9822 3049
rect 9644 2919 9678 2953
rect 9716 2919 9750 2953
rect 9788 2919 9822 2953
rect 9644 2823 9678 2857
rect 9716 2823 9750 2857
rect 9788 2823 9822 2857
rect 9644 2727 9678 2761
rect 9716 2727 9750 2761
rect 9788 2727 9822 2761
rect 9644 2631 9678 2665
rect 9716 2631 9750 2665
rect 9788 2631 9822 2665
rect 9644 2535 9678 2569
rect 9716 2535 9750 2569
rect 9788 2535 9822 2569
rect 9644 2439 9678 2473
rect 9716 2439 9750 2473
rect 9788 2439 9822 2473
rect 9644 2343 9678 2377
rect 9716 2343 9750 2377
rect 9788 2343 9822 2377
rect 9644 2247 9678 2281
rect 9716 2247 9750 2281
rect 9788 2247 9822 2281
rect 9644 2151 9678 2185
rect 9716 2151 9750 2185
rect 9788 2151 9822 2185
rect 9644 2055 9678 2089
rect 9716 2055 9750 2089
rect 9788 2055 9822 2089
rect 9644 1959 9678 1993
rect 9716 1959 9750 1993
rect 9788 1959 9822 1993
rect 9644 1863 9678 1897
rect 9716 1863 9750 1897
rect 9788 1863 9822 1897
rect 9644 1767 9678 1801
rect 9716 1767 9750 1801
rect 9788 1767 9822 1801
rect 9644 1671 9678 1705
rect 9716 1671 9750 1705
rect 9788 1671 9822 1705
rect 9644 1575 9678 1609
rect 9716 1575 9750 1609
rect 9788 1575 9822 1609
rect 9644 1479 9678 1513
rect 9716 1479 9750 1513
rect 9788 1479 9822 1513
rect 9644 1383 9678 1417
rect 9716 1383 9750 1417
rect 9788 1383 9822 1417
rect 9644 1287 9678 1321
rect 9716 1287 9750 1321
rect 9788 1287 9822 1321
rect 9644 1191 9678 1225
rect 9716 1191 9750 1225
rect 9788 1191 9822 1225
rect 9644 1095 9678 1129
rect 9716 1095 9750 1129
rect 9788 1095 9822 1129
rect 9644 999 9678 1033
rect 9716 999 9750 1033
rect 9788 999 9822 1033
rect 9644 903 9678 937
rect 9716 903 9750 937
rect 9788 903 9822 937
rect 9644 807 9678 841
rect 9716 807 9750 841
rect 9788 807 9822 841
rect 9644 711 9678 745
rect 9716 711 9750 745
rect 9788 711 9822 745
rect 9644 615 9678 649
rect 9716 615 9750 649
rect 9788 615 9822 649
rect 10056 3303 10090 3337
rect 10128 3303 10162 3337
rect 10200 3303 10234 3337
rect 10056 3207 10090 3241
rect 10128 3207 10162 3241
rect 10200 3207 10234 3241
rect 10056 3111 10090 3145
rect 10128 3111 10162 3145
rect 10200 3111 10234 3145
rect 10056 3015 10090 3049
rect 10128 3015 10162 3049
rect 10200 3015 10234 3049
rect 10056 2919 10090 2953
rect 10128 2919 10162 2953
rect 10200 2919 10234 2953
rect 10056 2823 10090 2857
rect 10128 2823 10162 2857
rect 10200 2823 10234 2857
rect 10056 2727 10090 2761
rect 10128 2727 10162 2761
rect 10200 2727 10234 2761
rect 10056 2631 10090 2665
rect 10128 2631 10162 2665
rect 10200 2631 10234 2665
rect 10056 2535 10090 2569
rect 10128 2535 10162 2569
rect 10200 2535 10234 2569
rect 10056 2439 10090 2473
rect 10128 2439 10162 2473
rect 10200 2439 10234 2473
rect 10056 2343 10090 2377
rect 10128 2343 10162 2377
rect 10200 2343 10234 2377
rect 10056 2247 10090 2281
rect 10128 2247 10162 2281
rect 10200 2247 10234 2281
rect 10056 2151 10090 2185
rect 10128 2151 10162 2185
rect 10200 2151 10234 2185
rect 10056 2055 10090 2089
rect 10128 2055 10162 2089
rect 10200 2055 10234 2089
rect 10056 1959 10090 1993
rect 10128 1959 10162 1993
rect 10200 1959 10234 1993
rect 10056 1863 10090 1897
rect 10128 1863 10162 1897
rect 10200 1863 10234 1897
rect 10056 1767 10090 1801
rect 10128 1767 10162 1801
rect 10200 1767 10234 1801
rect 10056 1671 10090 1705
rect 10128 1671 10162 1705
rect 10200 1671 10234 1705
rect 10056 1575 10090 1609
rect 10128 1575 10162 1609
rect 10200 1575 10234 1609
rect 10056 1479 10090 1513
rect 10128 1479 10162 1513
rect 10200 1479 10234 1513
rect 10056 1383 10090 1417
rect 10128 1383 10162 1417
rect 10200 1383 10234 1417
rect 10056 1287 10090 1321
rect 10128 1287 10162 1321
rect 10200 1287 10234 1321
rect 10056 1191 10090 1225
rect 10128 1191 10162 1225
rect 10200 1191 10234 1225
rect 10056 1095 10090 1129
rect 10128 1095 10162 1129
rect 10200 1095 10234 1129
rect 10056 999 10090 1033
rect 10128 999 10162 1033
rect 10200 999 10234 1033
rect 10056 903 10090 937
rect 10128 903 10162 937
rect 10200 903 10234 937
rect 10056 807 10090 841
rect 10128 807 10162 841
rect 10200 807 10234 841
rect 10056 711 10090 745
rect 10128 711 10162 745
rect 10200 711 10234 745
rect 10056 615 10090 649
rect 10128 615 10162 649
rect 10200 615 10234 649
rect 10468 3303 10502 3337
rect 10540 3303 10574 3337
rect 10612 3303 10646 3337
rect 10468 3207 10502 3241
rect 10540 3207 10574 3241
rect 10612 3207 10646 3241
rect 10468 3111 10502 3145
rect 10540 3111 10574 3145
rect 10612 3111 10646 3145
rect 10468 3015 10502 3049
rect 10540 3015 10574 3049
rect 10612 3015 10646 3049
rect 10468 2919 10502 2953
rect 10540 2919 10574 2953
rect 10612 2919 10646 2953
rect 10468 2823 10502 2857
rect 10540 2823 10574 2857
rect 10612 2823 10646 2857
rect 10468 2727 10502 2761
rect 10540 2727 10574 2761
rect 10612 2727 10646 2761
rect 10468 2631 10502 2665
rect 10540 2631 10574 2665
rect 10612 2631 10646 2665
rect 10468 2535 10502 2569
rect 10540 2535 10574 2569
rect 10612 2535 10646 2569
rect 10468 2439 10502 2473
rect 10540 2439 10574 2473
rect 10612 2439 10646 2473
rect 10468 2343 10502 2377
rect 10540 2343 10574 2377
rect 10612 2343 10646 2377
rect 10468 2247 10502 2281
rect 10540 2247 10574 2281
rect 10612 2247 10646 2281
rect 10468 2151 10502 2185
rect 10540 2151 10574 2185
rect 10612 2151 10646 2185
rect 10468 2055 10502 2089
rect 10540 2055 10574 2089
rect 10612 2055 10646 2089
rect 10468 1959 10502 1993
rect 10540 1959 10574 1993
rect 10612 1959 10646 1993
rect 10468 1863 10502 1897
rect 10540 1863 10574 1897
rect 10612 1863 10646 1897
rect 10468 1767 10502 1801
rect 10540 1767 10574 1801
rect 10612 1767 10646 1801
rect 10468 1671 10502 1705
rect 10540 1671 10574 1705
rect 10612 1671 10646 1705
rect 10468 1575 10502 1609
rect 10540 1575 10574 1609
rect 10612 1575 10646 1609
rect 10468 1479 10502 1513
rect 10540 1479 10574 1513
rect 10612 1479 10646 1513
rect 10468 1383 10502 1417
rect 10540 1383 10574 1417
rect 10612 1383 10646 1417
rect 10468 1287 10502 1321
rect 10540 1287 10574 1321
rect 10612 1287 10646 1321
rect 10468 1191 10502 1225
rect 10540 1191 10574 1225
rect 10612 1191 10646 1225
rect 10468 1095 10502 1129
rect 10540 1095 10574 1129
rect 10612 1095 10646 1129
rect 10468 999 10502 1033
rect 10540 999 10574 1033
rect 10612 999 10646 1033
rect 10468 903 10502 937
rect 10540 903 10574 937
rect 10612 903 10646 937
rect 10468 807 10502 841
rect 10540 807 10574 841
rect 10612 807 10646 841
rect 10468 711 10502 745
rect 10540 711 10574 745
rect 10612 711 10646 745
rect 10468 615 10502 649
rect 10540 615 10574 649
rect 10612 615 10646 649
rect 10880 3303 10914 3337
rect 10952 3303 10986 3337
rect 11024 3303 11058 3337
rect 10880 3207 10914 3241
rect 10952 3207 10986 3241
rect 11024 3207 11058 3241
rect 10880 3111 10914 3145
rect 10952 3111 10986 3145
rect 11024 3111 11058 3145
rect 10880 3015 10914 3049
rect 10952 3015 10986 3049
rect 11024 3015 11058 3049
rect 10880 2919 10914 2953
rect 10952 2919 10986 2953
rect 11024 2919 11058 2953
rect 10880 2823 10914 2857
rect 10952 2823 10986 2857
rect 11024 2823 11058 2857
rect 10880 2727 10914 2761
rect 10952 2727 10986 2761
rect 11024 2727 11058 2761
rect 10880 2631 10914 2665
rect 10952 2631 10986 2665
rect 11024 2631 11058 2665
rect 10880 2535 10914 2569
rect 10952 2535 10986 2569
rect 11024 2535 11058 2569
rect 10880 2439 10914 2473
rect 10952 2439 10986 2473
rect 11024 2439 11058 2473
rect 10880 2343 10914 2377
rect 10952 2343 10986 2377
rect 11024 2343 11058 2377
rect 10880 2247 10914 2281
rect 10952 2247 10986 2281
rect 11024 2247 11058 2281
rect 10880 2151 10914 2185
rect 10952 2151 10986 2185
rect 11024 2151 11058 2185
rect 10880 2055 10914 2089
rect 10952 2055 10986 2089
rect 11024 2055 11058 2089
rect 10880 1959 10914 1993
rect 10952 1959 10986 1993
rect 11024 1959 11058 1993
rect 10880 1863 10914 1897
rect 10952 1863 10986 1897
rect 11024 1863 11058 1897
rect 10880 1767 10914 1801
rect 10952 1767 10986 1801
rect 11024 1767 11058 1801
rect 10880 1671 10914 1705
rect 10952 1671 10986 1705
rect 11024 1671 11058 1705
rect 10880 1575 10914 1609
rect 10952 1575 10986 1609
rect 11024 1575 11058 1609
rect 10880 1479 10914 1513
rect 10952 1479 10986 1513
rect 11024 1479 11058 1513
rect 10880 1383 10914 1417
rect 10952 1383 10986 1417
rect 11024 1383 11058 1417
rect 10880 1287 10914 1321
rect 10952 1287 10986 1321
rect 11024 1287 11058 1321
rect 10880 1191 10914 1225
rect 10952 1191 10986 1225
rect 11024 1191 11058 1225
rect 10880 1095 10914 1129
rect 10952 1095 10986 1129
rect 11024 1095 11058 1129
rect 10880 999 10914 1033
rect 10952 999 10986 1033
rect 11024 999 11058 1033
rect 10880 903 10914 937
rect 10952 903 10986 937
rect 11024 903 11058 937
rect 10880 807 10914 841
rect 10952 807 10986 841
rect 11024 807 11058 841
rect 10880 711 10914 745
rect 10952 711 10986 745
rect 11024 711 11058 745
rect 10880 615 10914 649
rect 10952 615 10986 649
rect 11024 615 11058 649
rect 11328 3455 11331 3464
rect 11331 3455 11362 3464
rect 11328 3430 11362 3455
rect 11328 3387 11331 3392
rect 11331 3387 11362 3392
rect 11328 3358 11362 3387
rect 11328 3319 11331 3320
rect 11331 3319 11362 3320
rect 11328 3286 11362 3319
rect 11328 3217 11362 3248
rect 11328 3214 11331 3217
rect 11331 3214 11362 3217
rect 11328 3149 11362 3176
rect 11328 3142 11331 3149
rect 11331 3142 11362 3149
rect 11328 3081 11362 3104
rect 11328 3070 11331 3081
rect 11331 3070 11362 3081
rect 11328 3013 11362 3032
rect 11328 2998 11331 3013
rect 11331 2998 11362 3013
rect 11328 2945 11362 2960
rect 11328 2926 11331 2945
rect 11331 2926 11362 2945
rect 11328 2877 11362 2888
rect 11328 2854 11331 2877
rect 11331 2854 11362 2877
rect 11328 2809 11362 2816
rect 11328 2782 11331 2809
rect 11331 2782 11362 2809
rect 11328 2741 11362 2744
rect 11328 2710 11331 2741
rect 11331 2710 11362 2741
rect 11328 2639 11331 2672
rect 11331 2639 11362 2672
rect 11328 2638 11362 2639
rect 11328 2571 11331 2600
rect 11331 2571 11362 2600
rect 11328 2566 11362 2571
rect 11328 2503 11331 2528
rect 11331 2503 11362 2528
rect 11328 2494 11362 2503
rect 11328 2435 11331 2456
rect 11331 2435 11362 2456
rect 11328 2422 11362 2435
rect 11328 2367 11331 2384
rect 11331 2367 11362 2384
rect 11328 2350 11362 2367
rect 11328 2299 11331 2312
rect 11331 2299 11362 2312
rect 11328 2278 11362 2299
rect 11328 2231 11331 2240
rect 11331 2231 11362 2240
rect 11328 2206 11362 2231
rect 11328 2163 11331 2168
rect 11331 2163 11362 2168
rect 11328 2134 11362 2163
rect 11328 2095 11331 2096
rect 11331 2095 11362 2096
rect 11328 2062 11362 2095
rect 11328 1993 11362 2024
rect 11328 1990 11331 1993
rect 11331 1990 11362 1993
rect 11328 1925 11362 1952
rect 11328 1918 11331 1925
rect 11331 1918 11362 1925
rect 11328 1857 11362 1880
rect 11328 1846 11331 1857
rect 11331 1846 11362 1857
rect 11328 1789 11362 1808
rect 11328 1774 11331 1789
rect 11331 1774 11362 1789
rect 11328 1721 11362 1736
rect 11328 1702 11331 1721
rect 11331 1702 11362 1721
rect 11328 1653 11362 1664
rect 11328 1630 11331 1653
rect 11331 1630 11362 1653
rect 11328 1585 11362 1592
rect 11328 1558 11331 1585
rect 11331 1558 11362 1585
rect 11328 1517 11362 1520
rect 11328 1486 11331 1517
rect 11331 1486 11362 1517
rect 11328 1415 11331 1448
rect 11331 1415 11362 1448
rect 11328 1414 11362 1415
rect 11328 1347 11331 1376
rect 11331 1347 11362 1376
rect 11328 1342 11362 1347
rect 11328 1279 11331 1304
rect 11331 1279 11362 1304
rect 11328 1270 11362 1279
rect 11328 1211 11331 1232
rect 11331 1211 11362 1232
rect 11328 1198 11362 1211
rect 11328 1143 11331 1160
rect 11331 1143 11362 1160
rect 11328 1126 11362 1143
rect 11328 1075 11331 1088
rect 11331 1075 11362 1088
rect 11328 1054 11362 1075
rect 11328 1007 11331 1016
rect 11331 1007 11362 1016
rect 11328 982 11362 1007
rect 11328 939 11331 944
rect 11331 939 11362 944
rect 11328 910 11362 939
rect 11328 871 11331 872
rect 11331 871 11362 872
rect 11328 838 11362 871
rect 11328 769 11362 800
rect 11328 766 11331 769
rect 11331 766 11362 769
rect 11328 701 11362 728
rect 11328 694 11331 701
rect 11331 694 11362 701
rect 11328 633 11362 656
rect 11328 622 11331 633
rect 11331 622 11362 633
<< metal1 >>
rect 7157 3712 11389 3718
rect 7157 3684 7352 3712
rect 7386 3684 7501 3712
rect 7535 3684 7574 3712
rect 7608 3684 7646 3712
rect 7680 3684 7718 3712
rect 7752 3684 7790 3712
rect 7824 3684 7862 3712
rect 7896 3684 7934 3712
rect 7968 3684 8006 3712
rect 8040 3684 8078 3712
rect 8112 3684 8150 3712
rect 8184 3684 8222 3712
rect 8256 3684 8294 3712
rect 8328 3684 8366 3712
rect 8400 3684 8438 3712
rect 8472 3684 8510 3712
rect 8544 3684 8582 3712
rect 8616 3684 8654 3712
rect 8688 3684 8726 3712
rect 8760 3684 8798 3712
rect 8832 3684 8870 3712
rect 8904 3684 8942 3712
rect 8976 3684 9014 3712
rect 9048 3684 9086 3712
rect 9120 3684 9158 3712
rect 9192 3684 9230 3712
rect 9264 3684 9302 3712
rect 9336 3684 9374 3712
rect 9408 3684 9446 3712
rect 9480 3684 9518 3712
rect 9552 3684 9590 3712
rect 9624 3684 9662 3712
rect 9696 3684 9734 3712
rect 9768 3684 9806 3712
rect 9840 3684 9878 3712
rect 9912 3684 9950 3712
rect 9984 3684 10022 3712
rect 10056 3684 10094 3712
rect 10128 3684 10166 3712
rect 10200 3684 10238 3712
rect 10272 3684 10310 3712
rect 10344 3684 10382 3712
rect 10416 3684 10454 3712
rect 10488 3684 10526 3712
rect 10560 3684 10598 3712
rect 10632 3684 10670 3712
rect 10704 3684 10742 3712
rect 10776 3684 10814 3712
rect 10848 3684 10886 3712
rect 7157 3568 7220 3684
rect 10856 3678 10886 3684
rect 10920 3678 10958 3712
rect 10992 3678 11030 3712
rect 11064 3678 11102 3712
rect 11136 3678 11250 3712
rect 11284 3678 11389 3712
rect 10856 3568 11389 3678
rect 7157 3548 11389 3568
rect 7157 3514 7274 3548
rect 7308 3528 11328 3548
rect 7308 3514 7369 3528
tri 7369 3514 7383 3528 nw
tri 11273 3514 11287 3528 ne
rect 11287 3514 11328 3528
rect 11362 3514 11389 3548
rect 7157 3464 7335 3514
tri 7335 3480 7369 3514 nw
tri 11287 3494 11307 3514 ne
tri 7571 3464 7583 3476 se
rect 7583 3464 7763 3476
tri 7763 3464 7775 3476 sw
tri 7983 3464 7995 3476 se
rect 7995 3464 8175 3476
tri 8175 3464 8187 3476 sw
tri 8395 3464 8407 3476 se
rect 8407 3464 8587 3476
tri 8587 3464 8599 3476 sw
tri 8807 3464 8819 3476 se
rect 8819 3464 8999 3476
tri 8999 3464 9011 3476 sw
tri 9219 3464 9231 3476 se
rect 9231 3464 9411 3476
tri 9411 3464 9423 3476 sw
tri 9631 3464 9643 3476 se
rect 9643 3464 9823 3476
tri 9823 3464 9835 3476 sw
tri 10043 3464 10055 3476 se
rect 10055 3464 10235 3476
tri 10235 3464 10247 3476 sw
tri 10455 3464 10467 3476 se
rect 10467 3464 10647 3476
tri 10647 3464 10659 3476 sw
tri 10867 3464 10879 3476 se
rect 10879 3464 11059 3476
tri 11059 3464 11071 3476 sw
rect 11307 3464 11389 3514
rect 7157 3430 7274 3464
rect 7308 3430 7335 3464
tri 7537 3430 7571 3464 se
rect 7571 3430 7775 3464
tri 7775 3430 7809 3464 sw
tri 7949 3430 7983 3464 se
rect 7983 3430 8187 3464
tri 8187 3430 8221 3464 sw
tri 8361 3430 8395 3464 se
rect 8395 3430 8599 3464
tri 8599 3430 8633 3464 sw
tri 8773 3430 8807 3464 se
rect 8807 3430 9011 3464
tri 9011 3430 9045 3464 sw
tri 9185 3430 9219 3464 se
rect 9219 3430 9423 3464
tri 9423 3430 9457 3464 sw
tri 9597 3430 9631 3464 se
rect 9631 3430 9835 3464
tri 9835 3430 9869 3464 sw
tri 10009 3430 10043 3464 se
rect 10043 3430 10247 3464
tri 10247 3430 10281 3464 sw
tri 10421 3430 10455 3464 se
rect 10455 3430 10659 3464
tri 10659 3430 10693 3464 sw
tri 10833 3430 10867 3464 se
rect 10867 3430 11071 3464
tri 11071 3430 11105 3464 sw
rect 11307 3430 11328 3464
rect 11362 3430 11389 3464
rect 7157 3392 7335 3430
rect 7157 3358 7274 3392
rect 7308 3358 7335 3392
rect 7157 3320 7335 3358
rect 7157 3286 7274 3320
rect 7308 3286 7335 3320
rect 7157 3248 7335 3286
rect 7157 3214 7274 3248
rect 7308 3214 7335 3248
rect 7157 3176 7335 3214
rect 7157 3142 7274 3176
rect 7308 3142 7335 3176
rect 7157 3104 7335 3142
rect 7157 3070 7274 3104
rect 7308 3070 7335 3104
rect 7157 3032 7335 3070
rect 7157 2998 7274 3032
rect 7308 2998 7335 3032
rect 7157 2960 7335 2998
rect 7157 2926 7274 2960
rect 7308 2926 7335 2960
rect 7157 2888 7335 2926
rect 7157 2854 7274 2888
rect 7308 2854 7335 2888
rect 7157 2816 7335 2854
rect 7157 2782 7274 2816
rect 7308 2782 7335 2816
rect 7157 2744 7335 2782
rect 7157 2710 7274 2744
rect 7308 2710 7335 2744
rect 7157 2672 7335 2710
rect 7157 2638 7274 2672
rect 7308 2638 7335 2672
rect 7157 2600 7335 2638
rect 7157 2566 7274 2600
rect 7308 2566 7335 2600
rect 7157 2528 7335 2566
rect 7157 2494 7274 2528
rect 7308 2494 7335 2528
rect 7157 2456 7335 2494
rect 7157 2422 7274 2456
rect 7308 2422 7335 2456
rect 7157 2384 7335 2422
rect 7157 2350 7274 2384
rect 7308 2350 7335 2384
rect 7157 2312 7335 2350
rect 7157 2278 7274 2312
rect 7308 2278 7335 2312
rect 7157 2240 7335 2278
rect 7157 2206 7274 2240
rect 7308 2206 7335 2240
rect 7157 2168 7335 2206
rect 7157 2134 7274 2168
rect 7308 2134 7335 2168
rect 7157 2096 7335 2134
rect 7157 2062 7274 2096
rect 7308 2062 7335 2096
rect 7157 2024 7335 2062
rect 7157 1990 7274 2024
rect 7308 1990 7335 2024
rect 7157 1952 7335 1990
rect 7157 1918 7274 1952
rect 7308 1918 7335 1952
rect 7157 1880 7335 1918
rect 7157 1846 7274 1880
rect 7308 1846 7335 1880
rect 7157 1808 7335 1846
rect 7157 1774 7274 1808
rect 7308 1774 7335 1808
rect 7157 1736 7335 1774
rect 7157 1702 7274 1736
rect 7308 1702 7335 1736
rect 7157 1664 7335 1702
rect 7157 1630 7274 1664
rect 7308 1630 7335 1664
rect 7157 1592 7335 1630
rect 7157 1558 7274 1592
rect 7308 1558 7335 1592
rect 7157 1520 7335 1558
rect 7157 1486 7274 1520
rect 7308 1486 7335 1520
rect 7157 1448 7335 1486
rect 7157 1414 7274 1448
rect 7308 1414 7335 1448
rect 7157 1376 7335 1414
rect 7157 1342 7274 1376
rect 7308 1342 7335 1376
rect 7157 1304 7335 1342
rect 7157 1270 7274 1304
rect 7308 1270 7335 1304
rect 7157 1232 7335 1270
rect 7157 1198 7274 1232
rect 7308 1198 7335 1232
rect 7157 1160 7335 1198
rect 7157 1126 7274 1160
rect 7308 1126 7335 1160
rect 7157 1088 7335 1126
rect 7157 1054 7274 1088
rect 7308 1054 7335 1088
rect 7157 1016 7335 1054
rect 7157 982 7274 1016
rect 7308 982 7335 1016
rect 7157 944 7335 982
rect 7157 910 7274 944
rect 7308 910 7335 944
rect 7157 872 7335 910
rect 7157 838 7274 872
rect 7308 838 7335 872
rect 7157 800 7335 838
rect 7157 766 7274 800
rect 7308 766 7335 800
rect 7157 728 7335 766
rect 7157 694 7274 728
rect 7308 694 7335 728
rect 7157 656 7335 694
rect 7157 622 7274 656
rect 7308 622 7335 656
rect 7157 609 7335 622
tri 7523 3416 7537 3430 se
rect 7537 3416 7809 3430
tri 7809 3416 7823 3430 sw
rect 7523 3382 7823 3416
rect 7523 2050 7551 3382
rect 7795 2050 7823 3382
rect 7523 1993 7823 2050
rect 7523 1959 7584 1993
rect 7618 1959 7656 1993
rect 7690 1959 7728 1993
rect 7762 1959 7823 1993
rect 7523 1897 7823 1959
rect 7523 1863 7584 1897
rect 7618 1863 7656 1897
rect 7690 1863 7728 1897
rect 7762 1863 7823 1897
rect 7523 1801 7823 1863
rect 7523 1767 7584 1801
rect 7618 1767 7656 1801
rect 7690 1767 7728 1801
rect 7762 1767 7823 1801
rect 7523 1705 7823 1767
rect 7523 1671 7584 1705
rect 7618 1671 7656 1705
rect 7690 1671 7728 1705
rect 7762 1671 7823 1705
rect 7523 1609 7823 1671
rect 7523 1575 7584 1609
rect 7618 1575 7656 1609
rect 7690 1575 7728 1609
rect 7762 1575 7823 1609
rect 7523 1513 7823 1575
rect 7523 1479 7584 1513
rect 7618 1479 7656 1513
rect 7690 1479 7728 1513
rect 7762 1479 7823 1513
rect 7523 1417 7823 1479
rect 7523 1383 7584 1417
rect 7618 1383 7656 1417
rect 7690 1383 7728 1417
rect 7762 1383 7823 1417
rect 7523 1321 7823 1383
rect 7523 1287 7584 1321
rect 7618 1287 7656 1321
rect 7690 1287 7728 1321
rect 7762 1287 7823 1321
rect 7523 1225 7823 1287
rect 7523 1191 7584 1225
rect 7618 1191 7656 1225
rect 7690 1191 7728 1225
rect 7762 1191 7823 1225
rect 7523 1129 7823 1191
rect 7523 1095 7584 1129
rect 7618 1095 7656 1129
rect 7690 1095 7728 1129
rect 7762 1095 7823 1129
rect 7523 1033 7823 1095
rect 7523 999 7584 1033
rect 7618 999 7656 1033
rect 7690 999 7728 1033
rect 7762 999 7823 1033
rect 7523 937 7823 999
rect 7523 903 7584 937
rect 7618 903 7656 937
rect 7690 903 7728 937
rect 7762 903 7823 937
rect 7523 841 7823 903
rect 7523 807 7584 841
rect 7618 807 7656 841
rect 7690 807 7728 841
rect 7762 807 7823 841
rect 7523 745 7823 807
rect 7523 711 7584 745
rect 7618 711 7656 745
rect 7690 711 7728 745
rect 7762 711 7823 745
rect 7523 649 7823 711
rect 7523 615 7584 649
rect 7618 615 7656 649
rect 7690 615 7728 649
rect 7762 615 7823 649
rect 7523 536 7823 615
tri 7523 476 7583 536 ne
rect 7583 476 7763 536
tri 7763 476 7823 536 nw
tri 7935 3416 7949 3430 se
rect 7949 3416 8221 3430
tri 8221 3416 8235 3430 sw
rect 7935 3337 8235 3416
rect 7935 3303 7996 3337
rect 8030 3303 8068 3337
rect 8102 3303 8140 3337
rect 8174 3303 8235 3337
rect 7935 3241 8235 3303
rect 7935 3207 7996 3241
rect 8030 3207 8068 3241
rect 8102 3207 8140 3241
rect 8174 3207 8235 3241
rect 7935 3145 8235 3207
rect 7935 3111 7996 3145
rect 8030 3111 8068 3145
rect 8102 3111 8140 3145
rect 8174 3111 8235 3145
rect 7935 3049 8235 3111
rect 7935 3015 7996 3049
rect 8030 3015 8068 3049
rect 8102 3015 8140 3049
rect 8174 3015 8235 3049
rect 7935 2953 8235 3015
rect 7935 2919 7996 2953
rect 8030 2919 8068 2953
rect 8102 2919 8140 2953
rect 8174 2919 8235 2953
rect 7935 2857 8235 2919
rect 7935 2823 7996 2857
rect 8030 2823 8068 2857
rect 8102 2823 8140 2857
rect 8174 2823 8235 2857
rect 7935 2761 8235 2823
rect 7935 2727 7996 2761
rect 8030 2727 8068 2761
rect 8102 2727 8140 2761
rect 8174 2727 8235 2761
rect 7935 2665 8235 2727
rect 7935 2631 7996 2665
rect 8030 2631 8068 2665
rect 8102 2631 8140 2665
rect 8174 2631 8235 2665
rect 7935 2569 8235 2631
rect 7935 2535 7996 2569
rect 8030 2535 8068 2569
rect 8102 2535 8140 2569
rect 8174 2535 8235 2569
rect 7935 2473 8235 2535
rect 7935 2439 7996 2473
rect 8030 2439 8068 2473
rect 8102 2439 8140 2473
rect 8174 2439 8235 2473
rect 7935 2377 8235 2439
rect 7935 2343 7996 2377
rect 8030 2343 8068 2377
rect 8102 2343 8140 2377
rect 8174 2343 8235 2377
rect 7935 2281 8235 2343
rect 7935 2247 7996 2281
rect 8030 2247 8068 2281
rect 8102 2247 8140 2281
rect 8174 2247 8235 2281
rect 7935 2185 8235 2247
rect 7935 2151 7996 2185
rect 8030 2151 8068 2185
rect 8102 2151 8140 2185
rect 8174 2151 8235 2185
rect 7935 2089 8235 2151
rect 7935 2055 7996 2089
rect 8030 2055 8068 2089
rect 8102 2055 8140 2089
rect 8174 2055 8235 2089
rect 7935 1993 8235 2055
rect 7935 1959 7996 1993
rect 8030 1959 8068 1993
rect 8102 1959 8140 1993
rect 8174 1959 8235 1993
rect 7935 1897 8235 1959
rect 7935 1875 7996 1897
rect 8030 1875 8068 1897
rect 8102 1875 8140 1897
rect 8174 1875 8235 1897
tri 7793 316 7935 458 se
rect 7935 351 7963 1875
rect 8207 351 8235 1875
tri 8347 3416 8361 3430 se
rect 8361 3416 8633 3430
tri 8633 3416 8647 3430 sw
rect 8347 3382 8647 3416
rect 8347 2050 8375 3382
rect 8619 2050 8647 3382
rect 8347 1993 8647 2050
rect 8347 1959 8408 1993
rect 8442 1959 8480 1993
rect 8514 1959 8552 1993
rect 8586 1959 8647 1993
rect 8347 1897 8647 1959
rect 8347 1863 8408 1897
rect 8442 1863 8480 1897
rect 8514 1863 8552 1897
rect 8586 1863 8647 1897
rect 8347 1801 8647 1863
rect 8347 1767 8408 1801
rect 8442 1767 8480 1801
rect 8514 1767 8552 1801
rect 8586 1767 8647 1801
rect 8347 1705 8647 1767
rect 8347 1671 8408 1705
rect 8442 1671 8480 1705
rect 8514 1671 8552 1705
rect 8586 1671 8647 1705
rect 8347 1609 8647 1671
rect 8347 1575 8408 1609
rect 8442 1575 8480 1609
rect 8514 1575 8552 1609
rect 8586 1575 8647 1609
rect 8347 1513 8647 1575
rect 8347 1479 8408 1513
rect 8442 1479 8480 1513
rect 8514 1479 8552 1513
rect 8586 1479 8647 1513
rect 8347 1417 8647 1479
rect 8347 1383 8408 1417
rect 8442 1383 8480 1417
rect 8514 1383 8552 1417
rect 8586 1383 8647 1417
rect 8347 1321 8647 1383
rect 8347 1287 8408 1321
rect 8442 1287 8480 1321
rect 8514 1287 8552 1321
rect 8586 1287 8647 1321
rect 8347 1225 8647 1287
rect 8347 1191 8408 1225
rect 8442 1191 8480 1225
rect 8514 1191 8552 1225
rect 8586 1191 8647 1225
rect 8347 1129 8647 1191
rect 8347 1095 8408 1129
rect 8442 1095 8480 1129
rect 8514 1095 8552 1129
rect 8586 1095 8647 1129
rect 8347 1033 8647 1095
rect 8347 999 8408 1033
rect 8442 999 8480 1033
rect 8514 999 8552 1033
rect 8586 999 8647 1033
rect 8347 937 8647 999
rect 8347 903 8408 937
rect 8442 903 8480 937
rect 8514 903 8552 937
rect 8586 903 8647 937
rect 8347 841 8647 903
rect 8347 807 8408 841
rect 8442 807 8480 841
rect 8514 807 8552 841
rect 8586 807 8647 841
rect 8347 745 8647 807
rect 8347 711 8408 745
rect 8442 711 8480 745
rect 8514 711 8552 745
rect 8586 711 8647 745
rect 8347 649 8647 711
rect 8347 615 8408 649
rect 8442 615 8480 649
rect 8514 615 8552 649
rect 8586 615 8647 649
rect 8347 536 8647 615
tri 8347 476 8407 536 ne
rect 8407 476 8587 536
tri 8587 476 8647 536 nw
tri 8759 3416 8773 3430 se
rect 8773 3416 9045 3430
tri 9045 3416 9059 3430 sw
rect 8759 3337 9059 3416
rect 8759 3303 8820 3337
rect 8854 3303 8892 3337
rect 8926 3303 8964 3337
rect 8998 3303 9059 3337
rect 8759 3241 9059 3303
rect 8759 3207 8820 3241
rect 8854 3207 8892 3241
rect 8926 3207 8964 3241
rect 8998 3207 9059 3241
rect 8759 3145 9059 3207
rect 8759 3111 8820 3145
rect 8854 3111 8892 3145
rect 8926 3111 8964 3145
rect 8998 3111 9059 3145
rect 8759 3049 9059 3111
rect 8759 3015 8820 3049
rect 8854 3015 8892 3049
rect 8926 3015 8964 3049
rect 8998 3015 9059 3049
rect 8759 2953 9059 3015
rect 8759 2919 8820 2953
rect 8854 2919 8892 2953
rect 8926 2919 8964 2953
rect 8998 2919 9059 2953
rect 8759 2857 9059 2919
rect 8759 2823 8820 2857
rect 8854 2823 8892 2857
rect 8926 2823 8964 2857
rect 8998 2823 9059 2857
rect 8759 2761 9059 2823
rect 8759 2727 8820 2761
rect 8854 2727 8892 2761
rect 8926 2727 8964 2761
rect 8998 2727 9059 2761
rect 8759 2665 9059 2727
rect 8759 2631 8820 2665
rect 8854 2631 8892 2665
rect 8926 2631 8964 2665
rect 8998 2631 9059 2665
rect 8759 2569 9059 2631
rect 8759 2535 8820 2569
rect 8854 2535 8892 2569
rect 8926 2535 8964 2569
rect 8998 2535 9059 2569
rect 8759 2473 9059 2535
rect 8759 2439 8820 2473
rect 8854 2439 8892 2473
rect 8926 2439 8964 2473
rect 8998 2439 9059 2473
rect 8759 2377 9059 2439
rect 8759 2343 8820 2377
rect 8854 2343 8892 2377
rect 8926 2343 8964 2377
rect 8998 2343 9059 2377
rect 8759 2281 9059 2343
rect 8759 2247 8820 2281
rect 8854 2247 8892 2281
rect 8926 2247 8964 2281
rect 8998 2247 9059 2281
rect 8759 2185 9059 2247
rect 8759 2151 8820 2185
rect 8854 2151 8892 2185
rect 8926 2151 8964 2185
rect 8998 2151 9059 2185
rect 8759 2089 9059 2151
rect 8759 2055 8820 2089
rect 8854 2055 8892 2089
rect 8926 2055 8964 2089
rect 8998 2055 9059 2089
rect 8759 1993 9059 2055
rect 8759 1959 8820 1993
rect 8854 1959 8892 1993
rect 8926 1959 8964 1993
rect 8998 1959 9059 1993
rect 8759 1897 9059 1959
rect 8759 1875 8820 1897
rect 8854 1875 8892 1897
rect 8926 1875 8964 1897
rect 8998 1875 9059 1897
rect 7935 316 8235 351
tri 8235 316 8377 458 sw
tri 8617 316 8759 458 se
rect 8759 351 8787 1875
rect 9031 351 9059 1875
tri 9171 3416 9185 3430 se
rect 9185 3416 9457 3430
tri 9457 3416 9471 3430 sw
rect 9171 3382 9471 3416
rect 9171 2050 9199 3382
rect 9443 2050 9471 3382
rect 9171 1993 9471 2050
rect 9171 1959 9232 1993
rect 9266 1959 9304 1993
rect 9338 1959 9376 1993
rect 9410 1959 9471 1993
rect 9171 1897 9471 1959
rect 9171 1863 9232 1897
rect 9266 1863 9304 1897
rect 9338 1863 9376 1897
rect 9410 1863 9471 1897
rect 9171 1801 9471 1863
rect 9171 1767 9232 1801
rect 9266 1767 9304 1801
rect 9338 1767 9376 1801
rect 9410 1767 9471 1801
rect 9171 1705 9471 1767
rect 9171 1671 9232 1705
rect 9266 1671 9304 1705
rect 9338 1671 9376 1705
rect 9410 1671 9471 1705
rect 9171 1609 9471 1671
rect 9171 1575 9232 1609
rect 9266 1575 9304 1609
rect 9338 1575 9376 1609
rect 9410 1575 9471 1609
rect 9171 1513 9471 1575
rect 9171 1479 9232 1513
rect 9266 1479 9304 1513
rect 9338 1479 9376 1513
rect 9410 1479 9471 1513
rect 9171 1417 9471 1479
rect 9171 1383 9232 1417
rect 9266 1383 9304 1417
rect 9338 1383 9376 1417
rect 9410 1383 9471 1417
rect 9171 1321 9471 1383
rect 9171 1287 9232 1321
rect 9266 1287 9304 1321
rect 9338 1287 9376 1321
rect 9410 1287 9471 1321
rect 9171 1225 9471 1287
rect 9171 1191 9232 1225
rect 9266 1191 9304 1225
rect 9338 1191 9376 1225
rect 9410 1191 9471 1225
rect 9171 1129 9471 1191
rect 9171 1095 9232 1129
rect 9266 1095 9304 1129
rect 9338 1095 9376 1129
rect 9410 1095 9471 1129
rect 9171 1033 9471 1095
rect 9171 999 9232 1033
rect 9266 999 9304 1033
rect 9338 999 9376 1033
rect 9410 999 9471 1033
rect 9171 937 9471 999
rect 9171 903 9232 937
rect 9266 903 9304 937
rect 9338 903 9376 937
rect 9410 903 9471 937
rect 9171 841 9471 903
rect 9171 807 9232 841
rect 9266 807 9304 841
rect 9338 807 9376 841
rect 9410 807 9471 841
rect 9171 745 9471 807
rect 9171 711 9232 745
rect 9266 711 9304 745
rect 9338 711 9376 745
rect 9410 711 9471 745
rect 9171 649 9471 711
rect 9171 615 9232 649
rect 9266 615 9304 649
rect 9338 615 9376 649
rect 9410 615 9471 649
rect 9171 536 9471 615
tri 9171 476 9231 536 ne
rect 9231 476 9411 536
tri 9411 476 9471 536 nw
tri 9583 3416 9597 3430 se
rect 9597 3416 9869 3430
tri 9869 3416 9883 3430 sw
rect 9583 3337 9883 3416
rect 9583 3303 9644 3337
rect 9678 3303 9716 3337
rect 9750 3303 9788 3337
rect 9822 3303 9883 3337
rect 9583 3241 9883 3303
rect 9583 3207 9644 3241
rect 9678 3207 9716 3241
rect 9750 3207 9788 3241
rect 9822 3207 9883 3241
rect 9583 3145 9883 3207
rect 9583 3111 9644 3145
rect 9678 3111 9716 3145
rect 9750 3111 9788 3145
rect 9822 3111 9883 3145
rect 9583 3049 9883 3111
rect 9583 3015 9644 3049
rect 9678 3015 9716 3049
rect 9750 3015 9788 3049
rect 9822 3015 9883 3049
rect 9583 2953 9883 3015
rect 9583 2919 9644 2953
rect 9678 2919 9716 2953
rect 9750 2919 9788 2953
rect 9822 2919 9883 2953
rect 9583 2857 9883 2919
rect 9583 2823 9644 2857
rect 9678 2823 9716 2857
rect 9750 2823 9788 2857
rect 9822 2823 9883 2857
rect 9583 2761 9883 2823
rect 9583 2727 9644 2761
rect 9678 2727 9716 2761
rect 9750 2727 9788 2761
rect 9822 2727 9883 2761
rect 9583 2665 9883 2727
rect 9583 2631 9644 2665
rect 9678 2631 9716 2665
rect 9750 2631 9788 2665
rect 9822 2631 9883 2665
rect 9583 2569 9883 2631
rect 9583 2535 9644 2569
rect 9678 2535 9716 2569
rect 9750 2535 9788 2569
rect 9822 2535 9883 2569
rect 9583 2473 9883 2535
rect 9583 2439 9644 2473
rect 9678 2439 9716 2473
rect 9750 2439 9788 2473
rect 9822 2439 9883 2473
rect 9583 2377 9883 2439
rect 9583 2343 9644 2377
rect 9678 2343 9716 2377
rect 9750 2343 9788 2377
rect 9822 2343 9883 2377
rect 9583 2281 9883 2343
rect 9583 2247 9644 2281
rect 9678 2247 9716 2281
rect 9750 2247 9788 2281
rect 9822 2247 9883 2281
rect 9583 2185 9883 2247
rect 9583 2151 9644 2185
rect 9678 2151 9716 2185
rect 9750 2151 9788 2185
rect 9822 2151 9883 2185
rect 9583 2089 9883 2151
rect 9583 2055 9644 2089
rect 9678 2055 9716 2089
rect 9750 2055 9788 2089
rect 9822 2055 9883 2089
rect 9583 1993 9883 2055
rect 9583 1959 9644 1993
rect 9678 1959 9716 1993
rect 9750 1959 9788 1993
rect 9822 1959 9883 1993
rect 9583 1897 9883 1959
rect 9583 1875 9644 1897
rect 9678 1875 9716 1897
rect 9750 1875 9788 1897
rect 9822 1875 9883 1897
rect 8759 316 9059 351
tri 9059 316 9201 458 sw
tri 9441 316 9583 458 se
rect 9583 351 9611 1875
rect 9855 351 9883 1875
tri 9995 3416 10009 3430 se
rect 10009 3416 10281 3430
tri 10281 3416 10295 3430 sw
rect 9995 3382 10295 3416
rect 9995 2050 10023 3382
rect 10267 2050 10295 3382
rect 9995 1993 10295 2050
rect 9995 1959 10056 1993
rect 10090 1959 10128 1993
rect 10162 1959 10200 1993
rect 10234 1959 10295 1993
rect 9995 1897 10295 1959
rect 9995 1863 10056 1897
rect 10090 1863 10128 1897
rect 10162 1863 10200 1897
rect 10234 1863 10295 1897
rect 9995 1801 10295 1863
rect 9995 1767 10056 1801
rect 10090 1767 10128 1801
rect 10162 1767 10200 1801
rect 10234 1767 10295 1801
rect 9995 1705 10295 1767
rect 9995 1671 10056 1705
rect 10090 1671 10128 1705
rect 10162 1671 10200 1705
rect 10234 1671 10295 1705
rect 9995 1609 10295 1671
rect 9995 1575 10056 1609
rect 10090 1575 10128 1609
rect 10162 1575 10200 1609
rect 10234 1575 10295 1609
rect 9995 1513 10295 1575
rect 9995 1479 10056 1513
rect 10090 1479 10128 1513
rect 10162 1479 10200 1513
rect 10234 1479 10295 1513
rect 9995 1417 10295 1479
rect 9995 1383 10056 1417
rect 10090 1383 10128 1417
rect 10162 1383 10200 1417
rect 10234 1383 10295 1417
rect 9995 1321 10295 1383
rect 9995 1287 10056 1321
rect 10090 1287 10128 1321
rect 10162 1287 10200 1321
rect 10234 1287 10295 1321
rect 9995 1225 10295 1287
rect 9995 1191 10056 1225
rect 10090 1191 10128 1225
rect 10162 1191 10200 1225
rect 10234 1191 10295 1225
rect 9995 1129 10295 1191
rect 9995 1095 10056 1129
rect 10090 1095 10128 1129
rect 10162 1095 10200 1129
rect 10234 1095 10295 1129
rect 9995 1033 10295 1095
rect 9995 999 10056 1033
rect 10090 999 10128 1033
rect 10162 999 10200 1033
rect 10234 999 10295 1033
rect 9995 937 10295 999
rect 9995 903 10056 937
rect 10090 903 10128 937
rect 10162 903 10200 937
rect 10234 903 10295 937
rect 9995 841 10295 903
rect 9995 807 10056 841
rect 10090 807 10128 841
rect 10162 807 10200 841
rect 10234 807 10295 841
rect 9995 745 10295 807
rect 9995 711 10056 745
rect 10090 711 10128 745
rect 10162 711 10200 745
rect 10234 711 10295 745
rect 9995 649 10295 711
rect 9995 615 10056 649
rect 10090 615 10128 649
rect 10162 615 10200 649
rect 10234 615 10295 649
rect 9995 536 10295 615
tri 9995 476 10055 536 ne
rect 10055 476 10235 536
tri 10235 476 10295 536 nw
tri 10407 3416 10421 3430 se
rect 10421 3416 10693 3430
tri 10693 3416 10707 3430 sw
rect 10407 3337 10707 3416
rect 10407 3303 10468 3337
rect 10502 3303 10540 3337
rect 10574 3303 10612 3337
rect 10646 3303 10707 3337
rect 10407 3241 10707 3303
rect 10407 3207 10468 3241
rect 10502 3207 10540 3241
rect 10574 3207 10612 3241
rect 10646 3207 10707 3241
rect 10407 3145 10707 3207
rect 10407 3111 10468 3145
rect 10502 3111 10540 3145
rect 10574 3111 10612 3145
rect 10646 3111 10707 3145
rect 10407 3049 10707 3111
rect 10407 3015 10468 3049
rect 10502 3015 10540 3049
rect 10574 3015 10612 3049
rect 10646 3015 10707 3049
rect 10407 2953 10707 3015
rect 10407 2919 10468 2953
rect 10502 2919 10540 2953
rect 10574 2919 10612 2953
rect 10646 2919 10707 2953
rect 10407 2857 10707 2919
rect 10407 2823 10468 2857
rect 10502 2823 10540 2857
rect 10574 2823 10612 2857
rect 10646 2823 10707 2857
rect 10407 2761 10707 2823
rect 10407 2727 10468 2761
rect 10502 2727 10540 2761
rect 10574 2727 10612 2761
rect 10646 2727 10707 2761
rect 10407 2665 10707 2727
rect 10407 2631 10468 2665
rect 10502 2631 10540 2665
rect 10574 2631 10612 2665
rect 10646 2631 10707 2665
rect 10407 2569 10707 2631
rect 10407 2535 10468 2569
rect 10502 2535 10540 2569
rect 10574 2535 10612 2569
rect 10646 2535 10707 2569
rect 10407 2473 10707 2535
rect 10407 2439 10468 2473
rect 10502 2439 10540 2473
rect 10574 2439 10612 2473
rect 10646 2439 10707 2473
rect 10407 2377 10707 2439
rect 10407 2343 10468 2377
rect 10502 2343 10540 2377
rect 10574 2343 10612 2377
rect 10646 2343 10707 2377
rect 10407 2281 10707 2343
rect 10407 2247 10468 2281
rect 10502 2247 10540 2281
rect 10574 2247 10612 2281
rect 10646 2247 10707 2281
rect 10407 2185 10707 2247
rect 10407 2151 10468 2185
rect 10502 2151 10540 2185
rect 10574 2151 10612 2185
rect 10646 2151 10707 2185
rect 10407 2089 10707 2151
rect 10407 2055 10468 2089
rect 10502 2055 10540 2089
rect 10574 2055 10612 2089
rect 10646 2055 10707 2089
rect 10407 1993 10707 2055
rect 10407 1959 10468 1993
rect 10502 1959 10540 1993
rect 10574 1959 10612 1993
rect 10646 1959 10707 1993
rect 10407 1897 10707 1959
rect 10407 1875 10468 1897
rect 10502 1875 10540 1897
rect 10574 1875 10612 1897
rect 10646 1875 10707 1897
rect 9583 316 9883 351
tri 9883 316 10025 458 sw
tri 10265 316 10407 458 se
rect 10407 351 10435 1875
rect 10679 351 10707 1875
tri 10819 3416 10833 3430 se
rect 10833 3416 11105 3430
tri 11105 3416 11119 3430 sw
rect 10819 3382 11119 3416
rect 10819 2050 10847 3382
rect 11091 2050 11119 3382
rect 10819 1993 11119 2050
rect 10819 1959 10880 1993
rect 10914 1959 10952 1993
rect 10986 1959 11024 1993
rect 11058 1959 11119 1993
rect 10819 1897 11119 1959
rect 10819 1863 10880 1897
rect 10914 1863 10952 1897
rect 10986 1863 11024 1897
rect 11058 1863 11119 1897
rect 10819 1801 11119 1863
rect 10819 1767 10880 1801
rect 10914 1767 10952 1801
rect 10986 1767 11024 1801
rect 11058 1767 11119 1801
rect 10819 1705 11119 1767
rect 10819 1671 10880 1705
rect 10914 1671 10952 1705
rect 10986 1671 11024 1705
rect 11058 1671 11119 1705
rect 10819 1609 11119 1671
rect 10819 1575 10880 1609
rect 10914 1575 10952 1609
rect 10986 1575 11024 1609
rect 11058 1575 11119 1609
rect 10819 1513 11119 1575
rect 10819 1479 10880 1513
rect 10914 1479 10952 1513
rect 10986 1479 11024 1513
rect 11058 1479 11119 1513
rect 10819 1417 11119 1479
rect 10819 1383 10880 1417
rect 10914 1383 10952 1417
rect 10986 1383 11024 1417
rect 11058 1383 11119 1417
rect 10819 1321 11119 1383
rect 10819 1287 10880 1321
rect 10914 1287 10952 1321
rect 10986 1287 11024 1321
rect 11058 1287 11119 1321
rect 10819 1225 11119 1287
rect 10819 1191 10880 1225
rect 10914 1191 10952 1225
rect 10986 1191 11024 1225
rect 11058 1191 11119 1225
rect 10819 1129 11119 1191
rect 10819 1095 10880 1129
rect 10914 1095 10952 1129
rect 10986 1095 11024 1129
rect 11058 1095 11119 1129
rect 10819 1033 11119 1095
rect 10819 999 10880 1033
rect 10914 999 10952 1033
rect 10986 999 11024 1033
rect 11058 999 11119 1033
rect 10819 937 11119 999
rect 10819 903 10880 937
rect 10914 903 10952 937
rect 10986 903 11024 937
rect 11058 903 11119 937
rect 10819 841 11119 903
rect 10819 807 10880 841
rect 10914 807 10952 841
rect 10986 807 11024 841
rect 11058 807 11119 841
rect 10819 745 11119 807
rect 10819 711 10880 745
rect 10914 711 10952 745
rect 10986 711 11024 745
rect 11058 711 11119 745
rect 10819 649 11119 711
rect 10819 615 10880 649
rect 10914 615 10952 649
rect 10986 615 11024 649
rect 11058 615 11119 649
rect 10819 536 11119 615
rect 11307 3392 11389 3430
rect 11307 3358 11328 3392
rect 11362 3358 11389 3392
rect 11307 3320 11389 3358
rect 11307 3286 11328 3320
rect 11362 3286 11389 3320
rect 11307 3248 11389 3286
rect 11307 3214 11328 3248
rect 11362 3214 11389 3248
rect 11307 3176 11389 3214
rect 11307 3142 11328 3176
rect 11362 3142 11389 3176
rect 11307 3104 11389 3142
rect 11307 3070 11328 3104
rect 11362 3070 11389 3104
rect 11307 3032 11389 3070
rect 11307 2998 11328 3032
rect 11362 2998 11389 3032
rect 11307 2960 11389 2998
rect 11307 2926 11328 2960
rect 11362 2926 11389 2960
rect 11307 2888 11389 2926
rect 11307 2854 11328 2888
rect 11362 2854 11389 2888
rect 11307 2816 11389 2854
rect 11307 2782 11328 2816
rect 11362 2782 11389 2816
rect 11307 2744 11389 2782
rect 11307 2710 11328 2744
rect 11362 2710 11389 2744
rect 11307 2672 11389 2710
rect 11307 2638 11328 2672
rect 11362 2638 11389 2672
rect 11307 2600 11389 2638
rect 11307 2566 11328 2600
rect 11362 2566 11389 2600
rect 11307 2528 11389 2566
rect 11307 2494 11328 2528
rect 11362 2494 11389 2528
rect 11307 2456 11389 2494
rect 11307 2422 11328 2456
rect 11362 2422 11389 2456
rect 11307 2384 11389 2422
rect 11307 2350 11328 2384
rect 11362 2350 11389 2384
rect 11307 2312 11389 2350
rect 11307 2278 11328 2312
rect 11362 2278 11389 2312
rect 11307 2240 11389 2278
rect 11307 2206 11328 2240
rect 11362 2206 11389 2240
rect 11307 2168 11389 2206
rect 11307 2134 11328 2168
rect 11362 2134 11389 2168
rect 11307 2096 11389 2134
rect 11307 2062 11328 2096
rect 11362 2062 11389 2096
rect 11307 2024 11389 2062
rect 11307 1990 11328 2024
rect 11362 1990 11389 2024
rect 11307 1952 11389 1990
rect 11307 1918 11328 1952
rect 11362 1918 11389 1952
rect 11307 1880 11389 1918
rect 11307 1846 11328 1880
rect 11362 1846 11389 1880
rect 11307 1808 11389 1846
rect 11307 1774 11328 1808
rect 11362 1774 11389 1808
rect 11307 1736 11389 1774
rect 11307 1702 11328 1736
rect 11362 1702 11389 1736
rect 11307 1664 11389 1702
rect 11307 1630 11328 1664
rect 11362 1630 11389 1664
rect 11307 1592 11389 1630
rect 11307 1558 11328 1592
rect 11362 1558 11389 1592
rect 11307 1520 11389 1558
rect 11307 1486 11328 1520
rect 11362 1486 11389 1520
rect 11307 1448 11389 1486
rect 11307 1414 11328 1448
rect 11362 1414 11389 1448
rect 11307 1376 11389 1414
rect 11307 1342 11328 1376
rect 11362 1342 11389 1376
rect 11307 1304 11389 1342
rect 11307 1270 11328 1304
rect 11362 1270 11389 1304
rect 11307 1232 11389 1270
rect 11307 1198 11328 1232
rect 11362 1198 11389 1232
rect 11307 1160 11389 1198
rect 11307 1126 11328 1160
rect 11362 1126 11389 1160
rect 11307 1088 11389 1126
rect 11307 1054 11328 1088
rect 11362 1054 11389 1088
rect 11307 1016 11389 1054
rect 11307 982 11328 1016
rect 11362 982 11389 1016
rect 11307 944 11389 982
rect 11307 910 11328 944
rect 11362 910 11389 944
rect 11307 872 11389 910
rect 11307 838 11328 872
rect 11362 838 11389 872
rect 11307 800 11389 838
rect 11307 766 11328 800
rect 11362 766 11389 800
rect 11307 728 11389 766
rect 11307 694 11328 728
rect 11362 694 11389 728
rect 11307 656 11389 694
rect 11307 622 11328 656
rect 11362 622 11389 656
rect 11307 609 11389 622
tri 10819 476 10879 536 ne
rect 10879 476 11059 536
tri 11059 476 11119 536 nw
tri 11277 476 11307 506 se
rect 11307 476 11389 506
tri 11274 473 11277 476 se
rect 11277 473 11389 476
tri 11259 458 11274 473 se
rect 11274 458 11389 473
rect 10407 316 10707 351
tri 10707 316 10849 458 sw
tri 11117 316 11259 458 se
rect 11259 316 11389 458
rect 7157 288 11389 316
rect 7157 -20 7232 288
rect 10676 -20 11389 288
rect 7157 -48 11389 -20
<< via1 >>
rect 7220 3678 7352 3684
rect 7352 3678 7386 3684
rect 7386 3678 7501 3684
rect 7501 3678 7535 3684
rect 7535 3678 7574 3684
rect 7574 3678 7608 3684
rect 7608 3678 7646 3684
rect 7646 3678 7680 3684
rect 7680 3678 7718 3684
rect 7718 3678 7752 3684
rect 7752 3678 7790 3684
rect 7790 3678 7824 3684
rect 7824 3678 7862 3684
rect 7862 3678 7896 3684
rect 7896 3678 7934 3684
rect 7934 3678 7968 3684
rect 7968 3678 8006 3684
rect 8006 3678 8040 3684
rect 8040 3678 8078 3684
rect 8078 3678 8112 3684
rect 8112 3678 8150 3684
rect 8150 3678 8184 3684
rect 8184 3678 8222 3684
rect 8222 3678 8256 3684
rect 8256 3678 8294 3684
rect 8294 3678 8328 3684
rect 8328 3678 8366 3684
rect 8366 3678 8400 3684
rect 8400 3678 8438 3684
rect 8438 3678 8472 3684
rect 8472 3678 8510 3684
rect 8510 3678 8544 3684
rect 8544 3678 8582 3684
rect 8582 3678 8616 3684
rect 8616 3678 8654 3684
rect 8654 3678 8688 3684
rect 8688 3678 8726 3684
rect 8726 3678 8760 3684
rect 8760 3678 8798 3684
rect 8798 3678 8832 3684
rect 8832 3678 8870 3684
rect 8870 3678 8904 3684
rect 8904 3678 8942 3684
rect 8942 3678 8976 3684
rect 8976 3678 9014 3684
rect 9014 3678 9048 3684
rect 9048 3678 9086 3684
rect 9086 3678 9120 3684
rect 9120 3678 9158 3684
rect 9158 3678 9192 3684
rect 9192 3678 9230 3684
rect 9230 3678 9264 3684
rect 9264 3678 9302 3684
rect 9302 3678 9336 3684
rect 9336 3678 9374 3684
rect 9374 3678 9408 3684
rect 9408 3678 9446 3684
rect 9446 3678 9480 3684
rect 9480 3678 9518 3684
rect 9518 3678 9552 3684
rect 9552 3678 9590 3684
rect 9590 3678 9624 3684
rect 9624 3678 9662 3684
rect 9662 3678 9696 3684
rect 9696 3678 9734 3684
rect 9734 3678 9768 3684
rect 9768 3678 9806 3684
rect 9806 3678 9840 3684
rect 9840 3678 9878 3684
rect 9878 3678 9912 3684
rect 9912 3678 9950 3684
rect 9950 3678 9984 3684
rect 9984 3678 10022 3684
rect 10022 3678 10056 3684
rect 10056 3678 10094 3684
rect 10094 3678 10128 3684
rect 10128 3678 10166 3684
rect 10166 3678 10200 3684
rect 10200 3678 10238 3684
rect 10238 3678 10272 3684
rect 10272 3678 10310 3684
rect 10310 3678 10344 3684
rect 10344 3678 10382 3684
rect 10382 3678 10416 3684
rect 10416 3678 10454 3684
rect 10454 3678 10488 3684
rect 10488 3678 10526 3684
rect 10526 3678 10560 3684
rect 10560 3678 10598 3684
rect 10598 3678 10632 3684
rect 10632 3678 10670 3684
rect 10670 3678 10704 3684
rect 10704 3678 10742 3684
rect 10742 3678 10776 3684
rect 10776 3678 10814 3684
rect 10814 3678 10848 3684
rect 10848 3678 10856 3684
rect 7220 3568 10856 3678
rect 7551 3337 7795 3382
rect 7551 3303 7584 3337
rect 7584 3303 7618 3337
rect 7618 3303 7656 3337
rect 7656 3303 7690 3337
rect 7690 3303 7728 3337
rect 7728 3303 7762 3337
rect 7762 3303 7795 3337
rect 7551 3241 7795 3303
rect 7551 3207 7584 3241
rect 7584 3207 7618 3241
rect 7618 3207 7656 3241
rect 7656 3207 7690 3241
rect 7690 3207 7728 3241
rect 7728 3207 7762 3241
rect 7762 3207 7795 3241
rect 7551 3145 7795 3207
rect 7551 3111 7584 3145
rect 7584 3111 7618 3145
rect 7618 3111 7656 3145
rect 7656 3111 7690 3145
rect 7690 3111 7728 3145
rect 7728 3111 7762 3145
rect 7762 3111 7795 3145
rect 7551 3049 7795 3111
rect 7551 3015 7584 3049
rect 7584 3015 7618 3049
rect 7618 3015 7656 3049
rect 7656 3015 7690 3049
rect 7690 3015 7728 3049
rect 7728 3015 7762 3049
rect 7762 3015 7795 3049
rect 7551 2953 7795 3015
rect 7551 2919 7584 2953
rect 7584 2919 7618 2953
rect 7618 2919 7656 2953
rect 7656 2919 7690 2953
rect 7690 2919 7728 2953
rect 7728 2919 7762 2953
rect 7762 2919 7795 2953
rect 7551 2857 7795 2919
rect 7551 2823 7584 2857
rect 7584 2823 7618 2857
rect 7618 2823 7656 2857
rect 7656 2823 7690 2857
rect 7690 2823 7728 2857
rect 7728 2823 7762 2857
rect 7762 2823 7795 2857
rect 7551 2761 7795 2823
rect 7551 2727 7584 2761
rect 7584 2727 7618 2761
rect 7618 2727 7656 2761
rect 7656 2727 7690 2761
rect 7690 2727 7728 2761
rect 7728 2727 7762 2761
rect 7762 2727 7795 2761
rect 7551 2665 7795 2727
rect 7551 2631 7584 2665
rect 7584 2631 7618 2665
rect 7618 2631 7656 2665
rect 7656 2631 7690 2665
rect 7690 2631 7728 2665
rect 7728 2631 7762 2665
rect 7762 2631 7795 2665
rect 7551 2569 7795 2631
rect 7551 2535 7584 2569
rect 7584 2535 7618 2569
rect 7618 2535 7656 2569
rect 7656 2535 7690 2569
rect 7690 2535 7728 2569
rect 7728 2535 7762 2569
rect 7762 2535 7795 2569
rect 7551 2473 7795 2535
rect 7551 2439 7584 2473
rect 7584 2439 7618 2473
rect 7618 2439 7656 2473
rect 7656 2439 7690 2473
rect 7690 2439 7728 2473
rect 7728 2439 7762 2473
rect 7762 2439 7795 2473
rect 7551 2377 7795 2439
rect 7551 2343 7584 2377
rect 7584 2343 7618 2377
rect 7618 2343 7656 2377
rect 7656 2343 7690 2377
rect 7690 2343 7728 2377
rect 7728 2343 7762 2377
rect 7762 2343 7795 2377
rect 7551 2281 7795 2343
rect 7551 2247 7584 2281
rect 7584 2247 7618 2281
rect 7618 2247 7656 2281
rect 7656 2247 7690 2281
rect 7690 2247 7728 2281
rect 7728 2247 7762 2281
rect 7762 2247 7795 2281
rect 7551 2185 7795 2247
rect 7551 2151 7584 2185
rect 7584 2151 7618 2185
rect 7618 2151 7656 2185
rect 7656 2151 7690 2185
rect 7690 2151 7728 2185
rect 7728 2151 7762 2185
rect 7762 2151 7795 2185
rect 7551 2089 7795 2151
rect 7551 2055 7584 2089
rect 7584 2055 7618 2089
rect 7618 2055 7656 2089
rect 7656 2055 7690 2089
rect 7690 2055 7728 2089
rect 7728 2055 7762 2089
rect 7762 2055 7795 2089
rect 7551 2050 7795 2055
rect 7963 1863 7996 1875
rect 7996 1863 8030 1875
rect 8030 1863 8068 1875
rect 8068 1863 8102 1875
rect 8102 1863 8140 1875
rect 8140 1863 8174 1875
rect 8174 1863 8207 1875
rect 7963 1801 8207 1863
rect 7963 1767 7996 1801
rect 7996 1767 8030 1801
rect 8030 1767 8068 1801
rect 8068 1767 8102 1801
rect 8102 1767 8140 1801
rect 8140 1767 8174 1801
rect 8174 1767 8207 1801
rect 7963 1705 8207 1767
rect 7963 1671 7996 1705
rect 7996 1671 8030 1705
rect 8030 1671 8068 1705
rect 8068 1671 8102 1705
rect 8102 1671 8140 1705
rect 8140 1671 8174 1705
rect 8174 1671 8207 1705
rect 7963 1609 8207 1671
rect 7963 1575 7996 1609
rect 7996 1575 8030 1609
rect 8030 1575 8068 1609
rect 8068 1575 8102 1609
rect 8102 1575 8140 1609
rect 8140 1575 8174 1609
rect 8174 1575 8207 1609
rect 7963 1513 8207 1575
rect 7963 1479 7996 1513
rect 7996 1479 8030 1513
rect 8030 1479 8068 1513
rect 8068 1479 8102 1513
rect 8102 1479 8140 1513
rect 8140 1479 8174 1513
rect 8174 1479 8207 1513
rect 7963 1417 8207 1479
rect 7963 1383 7996 1417
rect 7996 1383 8030 1417
rect 8030 1383 8068 1417
rect 8068 1383 8102 1417
rect 8102 1383 8140 1417
rect 8140 1383 8174 1417
rect 8174 1383 8207 1417
rect 7963 1321 8207 1383
rect 7963 1287 7996 1321
rect 7996 1287 8030 1321
rect 8030 1287 8068 1321
rect 8068 1287 8102 1321
rect 8102 1287 8140 1321
rect 8140 1287 8174 1321
rect 8174 1287 8207 1321
rect 7963 1225 8207 1287
rect 7963 1191 7996 1225
rect 7996 1191 8030 1225
rect 8030 1191 8068 1225
rect 8068 1191 8102 1225
rect 8102 1191 8140 1225
rect 8140 1191 8174 1225
rect 8174 1191 8207 1225
rect 7963 1129 8207 1191
rect 7963 1095 7996 1129
rect 7996 1095 8030 1129
rect 8030 1095 8068 1129
rect 8068 1095 8102 1129
rect 8102 1095 8140 1129
rect 8140 1095 8174 1129
rect 8174 1095 8207 1129
rect 7963 1033 8207 1095
rect 7963 999 7996 1033
rect 7996 999 8030 1033
rect 8030 999 8068 1033
rect 8068 999 8102 1033
rect 8102 999 8140 1033
rect 8140 999 8174 1033
rect 8174 999 8207 1033
rect 7963 937 8207 999
rect 7963 903 7996 937
rect 7996 903 8030 937
rect 8030 903 8068 937
rect 8068 903 8102 937
rect 8102 903 8140 937
rect 8140 903 8174 937
rect 8174 903 8207 937
rect 7963 841 8207 903
rect 7963 807 7996 841
rect 7996 807 8030 841
rect 8030 807 8068 841
rect 8068 807 8102 841
rect 8102 807 8140 841
rect 8140 807 8174 841
rect 8174 807 8207 841
rect 7963 745 8207 807
rect 7963 711 7996 745
rect 7996 711 8030 745
rect 8030 711 8068 745
rect 8068 711 8102 745
rect 8102 711 8140 745
rect 8140 711 8174 745
rect 8174 711 8207 745
rect 7963 649 8207 711
rect 7963 615 7996 649
rect 7996 615 8030 649
rect 8030 615 8068 649
rect 8068 615 8102 649
rect 8102 615 8140 649
rect 8140 615 8174 649
rect 8174 615 8207 649
rect 7963 351 8207 615
rect 8375 3337 8619 3382
rect 8375 3303 8408 3337
rect 8408 3303 8442 3337
rect 8442 3303 8480 3337
rect 8480 3303 8514 3337
rect 8514 3303 8552 3337
rect 8552 3303 8586 3337
rect 8586 3303 8619 3337
rect 8375 3241 8619 3303
rect 8375 3207 8408 3241
rect 8408 3207 8442 3241
rect 8442 3207 8480 3241
rect 8480 3207 8514 3241
rect 8514 3207 8552 3241
rect 8552 3207 8586 3241
rect 8586 3207 8619 3241
rect 8375 3145 8619 3207
rect 8375 3111 8408 3145
rect 8408 3111 8442 3145
rect 8442 3111 8480 3145
rect 8480 3111 8514 3145
rect 8514 3111 8552 3145
rect 8552 3111 8586 3145
rect 8586 3111 8619 3145
rect 8375 3049 8619 3111
rect 8375 3015 8408 3049
rect 8408 3015 8442 3049
rect 8442 3015 8480 3049
rect 8480 3015 8514 3049
rect 8514 3015 8552 3049
rect 8552 3015 8586 3049
rect 8586 3015 8619 3049
rect 8375 2953 8619 3015
rect 8375 2919 8408 2953
rect 8408 2919 8442 2953
rect 8442 2919 8480 2953
rect 8480 2919 8514 2953
rect 8514 2919 8552 2953
rect 8552 2919 8586 2953
rect 8586 2919 8619 2953
rect 8375 2857 8619 2919
rect 8375 2823 8408 2857
rect 8408 2823 8442 2857
rect 8442 2823 8480 2857
rect 8480 2823 8514 2857
rect 8514 2823 8552 2857
rect 8552 2823 8586 2857
rect 8586 2823 8619 2857
rect 8375 2761 8619 2823
rect 8375 2727 8408 2761
rect 8408 2727 8442 2761
rect 8442 2727 8480 2761
rect 8480 2727 8514 2761
rect 8514 2727 8552 2761
rect 8552 2727 8586 2761
rect 8586 2727 8619 2761
rect 8375 2665 8619 2727
rect 8375 2631 8408 2665
rect 8408 2631 8442 2665
rect 8442 2631 8480 2665
rect 8480 2631 8514 2665
rect 8514 2631 8552 2665
rect 8552 2631 8586 2665
rect 8586 2631 8619 2665
rect 8375 2569 8619 2631
rect 8375 2535 8408 2569
rect 8408 2535 8442 2569
rect 8442 2535 8480 2569
rect 8480 2535 8514 2569
rect 8514 2535 8552 2569
rect 8552 2535 8586 2569
rect 8586 2535 8619 2569
rect 8375 2473 8619 2535
rect 8375 2439 8408 2473
rect 8408 2439 8442 2473
rect 8442 2439 8480 2473
rect 8480 2439 8514 2473
rect 8514 2439 8552 2473
rect 8552 2439 8586 2473
rect 8586 2439 8619 2473
rect 8375 2377 8619 2439
rect 8375 2343 8408 2377
rect 8408 2343 8442 2377
rect 8442 2343 8480 2377
rect 8480 2343 8514 2377
rect 8514 2343 8552 2377
rect 8552 2343 8586 2377
rect 8586 2343 8619 2377
rect 8375 2281 8619 2343
rect 8375 2247 8408 2281
rect 8408 2247 8442 2281
rect 8442 2247 8480 2281
rect 8480 2247 8514 2281
rect 8514 2247 8552 2281
rect 8552 2247 8586 2281
rect 8586 2247 8619 2281
rect 8375 2185 8619 2247
rect 8375 2151 8408 2185
rect 8408 2151 8442 2185
rect 8442 2151 8480 2185
rect 8480 2151 8514 2185
rect 8514 2151 8552 2185
rect 8552 2151 8586 2185
rect 8586 2151 8619 2185
rect 8375 2089 8619 2151
rect 8375 2055 8408 2089
rect 8408 2055 8442 2089
rect 8442 2055 8480 2089
rect 8480 2055 8514 2089
rect 8514 2055 8552 2089
rect 8552 2055 8586 2089
rect 8586 2055 8619 2089
rect 8375 2050 8619 2055
rect 8787 1863 8820 1875
rect 8820 1863 8854 1875
rect 8854 1863 8892 1875
rect 8892 1863 8926 1875
rect 8926 1863 8964 1875
rect 8964 1863 8998 1875
rect 8998 1863 9031 1875
rect 8787 1801 9031 1863
rect 8787 1767 8820 1801
rect 8820 1767 8854 1801
rect 8854 1767 8892 1801
rect 8892 1767 8926 1801
rect 8926 1767 8964 1801
rect 8964 1767 8998 1801
rect 8998 1767 9031 1801
rect 8787 1705 9031 1767
rect 8787 1671 8820 1705
rect 8820 1671 8854 1705
rect 8854 1671 8892 1705
rect 8892 1671 8926 1705
rect 8926 1671 8964 1705
rect 8964 1671 8998 1705
rect 8998 1671 9031 1705
rect 8787 1609 9031 1671
rect 8787 1575 8820 1609
rect 8820 1575 8854 1609
rect 8854 1575 8892 1609
rect 8892 1575 8926 1609
rect 8926 1575 8964 1609
rect 8964 1575 8998 1609
rect 8998 1575 9031 1609
rect 8787 1513 9031 1575
rect 8787 1479 8820 1513
rect 8820 1479 8854 1513
rect 8854 1479 8892 1513
rect 8892 1479 8926 1513
rect 8926 1479 8964 1513
rect 8964 1479 8998 1513
rect 8998 1479 9031 1513
rect 8787 1417 9031 1479
rect 8787 1383 8820 1417
rect 8820 1383 8854 1417
rect 8854 1383 8892 1417
rect 8892 1383 8926 1417
rect 8926 1383 8964 1417
rect 8964 1383 8998 1417
rect 8998 1383 9031 1417
rect 8787 1321 9031 1383
rect 8787 1287 8820 1321
rect 8820 1287 8854 1321
rect 8854 1287 8892 1321
rect 8892 1287 8926 1321
rect 8926 1287 8964 1321
rect 8964 1287 8998 1321
rect 8998 1287 9031 1321
rect 8787 1225 9031 1287
rect 8787 1191 8820 1225
rect 8820 1191 8854 1225
rect 8854 1191 8892 1225
rect 8892 1191 8926 1225
rect 8926 1191 8964 1225
rect 8964 1191 8998 1225
rect 8998 1191 9031 1225
rect 8787 1129 9031 1191
rect 8787 1095 8820 1129
rect 8820 1095 8854 1129
rect 8854 1095 8892 1129
rect 8892 1095 8926 1129
rect 8926 1095 8964 1129
rect 8964 1095 8998 1129
rect 8998 1095 9031 1129
rect 8787 1033 9031 1095
rect 8787 999 8820 1033
rect 8820 999 8854 1033
rect 8854 999 8892 1033
rect 8892 999 8926 1033
rect 8926 999 8964 1033
rect 8964 999 8998 1033
rect 8998 999 9031 1033
rect 8787 937 9031 999
rect 8787 903 8820 937
rect 8820 903 8854 937
rect 8854 903 8892 937
rect 8892 903 8926 937
rect 8926 903 8964 937
rect 8964 903 8998 937
rect 8998 903 9031 937
rect 8787 841 9031 903
rect 8787 807 8820 841
rect 8820 807 8854 841
rect 8854 807 8892 841
rect 8892 807 8926 841
rect 8926 807 8964 841
rect 8964 807 8998 841
rect 8998 807 9031 841
rect 8787 745 9031 807
rect 8787 711 8820 745
rect 8820 711 8854 745
rect 8854 711 8892 745
rect 8892 711 8926 745
rect 8926 711 8964 745
rect 8964 711 8998 745
rect 8998 711 9031 745
rect 8787 649 9031 711
rect 8787 615 8820 649
rect 8820 615 8854 649
rect 8854 615 8892 649
rect 8892 615 8926 649
rect 8926 615 8964 649
rect 8964 615 8998 649
rect 8998 615 9031 649
rect 8787 351 9031 615
rect 9199 3337 9443 3382
rect 9199 3303 9232 3337
rect 9232 3303 9266 3337
rect 9266 3303 9304 3337
rect 9304 3303 9338 3337
rect 9338 3303 9376 3337
rect 9376 3303 9410 3337
rect 9410 3303 9443 3337
rect 9199 3241 9443 3303
rect 9199 3207 9232 3241
rect 9232 3207 9266 3241
rect 9266 3207 9304 3241
rect 9304 3207 9338 3241
rect 9338 3207 9376 3241
rect 9376 3207 9410 3241
rect 9410 3207 9443 3241
rect 9199 3145 9443 3207
rect 9199 3111 9232 3145
rect 9232 3111 9266 3145
rect 9266 3111 9304 3145
rect 9304 3111 9338 3145
rect 9338 3111 9376 3145
rect 9376 3111 9410 3145
rect 9410 3111 9443 3145
rect 9199 3049 9443 3111
rect 9199 3015 9232 3049
rect 9232 3015 9266 3049
rect 9266 3015 9304 3049
rect 9304 3015 9338 3049
rect 9338 3015 9376 3049
rect 9376 3015 9410 3049
rect 9410 3015 9443 3049
rect 9199 2953 9443 3015
rect 9199 2919 9232 2953
rect 9232 2919 9266 2953
rect 9266 2919 9304 2953
rect 9304 2919 9338 2953
rect 9338 2919 9376 2953
rect 9376 2919 9410 2953
rect 9410 2919 9443 2953
rect 9199 2857 9443 2919
rect 9199 2823 9232 2857
rect 9232 2823 9266 2857
rect 9266 2823 9304 2857
rect 9304 2823 9338 2857
rect 9338 2823 9376 2857
rect 9376 2823 9410 2857
rect 9410 2823 9443 2857
rect 9199 2761 9443 2823
rect 9199 2727 9232 2761
rect 9232 2727 9266 2761
rect 9266 2727 9304 2761
rect 9304 2727 9338 2761
rect 9338 2727 9376 2761
rect 9376 2727 9410 2761
rect 9410 2727 9443 2761
rect 9199 2665 9443 2727
rect 9199 2631 9232 2665
rect 9232 2631 9266 2665
rect 9266 2631 9304 2665
rect 9304 2631 9338 2665
rect 9338 2631 9376 2665
rect 9376 2631 9410 2665
rect 9410 2631 9443 2665
rect 9199 2569 9443 2631
rect 9199 2535 9232 2569
rect 9232 2535 9266 2569
rect 9266 2535 9304 2569
rect 9304 2535 9338 2569
rect 9338 2535 9376 2569
rect 9376 2535 9410 2569
rect 9410 2535 9443 2569
rect 9199 2473 9443 2535
rect 9199 2439 9232 2473
rect 9232 2439 9266 2473
rect 9266 2439 9304 2473
rect 9304 2439 9338 2473
rect 9338 2439 9376 2473
rect 9376 2439 9410 2473
rect 9410 2439 9443 2473
rect 9199 2377 9443 2439
rect 9199 2343 9232 2377
rect 9232 2343 9266 2377
rect 9266 2343 9304 2377
rect 9304 2343 9338 2377
rect 9338 2343 9376 2377
rect 9376 2343 9410 2377
rect 9410 2343 9443 2377
rect 9199 2281 9443 2343
rect 9199 2247 9232 2281
rect 9232 2247 9266 2281
rect 9266 2247 9304 2281
rect 9304 2247 9338 2281
rect 9338 2247 9376 2281
rect 9376 2247 9410 2281
rect 9410 2247 9443 2281
rect 9199 2185 9443 2247
rect 9199 2151 9232 2185
rect 9232 2151 9266 2185
rect 9266 2151 9304 2185
rect 9304 2151 9338 2185
rect 9338 2151 9376 2185
rect 9376 2151 9410 2185
rect 9410 2151 9443 2185
rect 9199 2089 9443 2151
rect 9199 2055 9232 2089
rect 9232 2055 9266 2089
rect 9266 2055 9304 2089
rect 9304 2055 9338 2089
rect 9338 2055 9376 2089
rect 9376 2055 9410 2089
rect 9410 2055 9443 2089
rect 9199 2050 9443 2055
rect 9611 1863 9644 1875
rect 9644 1863 9678 1875
rect 9678 1863 9716 1875
rect 9716 1863 9750 1875
rect 9750 1863 9788 1875
rect 9788 1863 9822 1875
rect 9822 1863 9855 1875
rect 9611 1801 9855 1863
rect 9611 1767 9644 1801
rect 9644 1767 9678 1801
rect 9678 1767 9716 1801
rect 9716 1767 9750 1801
rect 9750 1767 9788 1801
rect 9788 1767 9822 1801
rect 9822 1767 9855 1801
rect 9611 1705 9855 1767
rect 9611 1671 9644 1705
rect 9644 1671 9678 1705
rect 9678 1671 9716 1705
rect 9716 1671 9750 1705
rect 9750 1671 9788 1705
rect 9788 1671 9822 1705
rect 9822 1671 9855 1705
rect 9611 1609 9855 1671
rect 9611 1575 9644 1609
rect 9644 1575 9678 1609
rect 9678 1575 9716 1609
rect 9716 1575 9750 1609
rect 9750 1575 9788 1609
rect 9788 1575 9822 1609
rect 9822 1575 9855 1609
rect 9611 1513 9855 1575
rect 9611 1479 9644 1513
rect 9644 1479 9678 1513
rect 9678 1479 9716 1513
rect 9716 1479 9750 1513
rect 9750 1479 9788 1513
rect 9788 1479 9822 1513
rect 9822 1479 9855 1513
rect 9611 1417 9855 1479
rect 9611 1383 9644 1417
rect 9644 1383 9678 1417
rect 9678 1383 9716 1417
rect 9716 1383 9750 1417
rect 9750 1383 9788 1417
rect 9788 1383 9822 1417
rect 9822 1383 9855 1417
rect 9611 1321 9855 1383
rect 9611 1287 9644 1321
rect 9644 1287 9678 1321
rect 9678 1287 9716 1321
rect 9716 1287 9750 1321
rect 9750 1287 9788 1321
rect 9788 1287 9822 1321
rect 9822 1287 9855 1321
rect 9611 1225 9855 1287
rect 9611 1191 9644 1225
rect 9644 1191 9678 1225
rect 9678 1191 9716 1225
rect 9716 1191 9750 1225
rect 9750 1191 9788 1225
rect 9788 1191 9822 1225
rect 9822 1191 9855 1225
rect 9611 1129 9855 1191
rect 9611 1095 9644 1129
rect 9644 1095 9678 1129
rect 9678 1095 9716 1129
rect 9716 1095 9750 1129
rect 9750 1095 9788 1129
rect 9788 1095 9822 1129
rect 9822 1095 9855 1129
rect 9611 1033 9855 1095
rect 9611 999 9644 1033
rect 9644 999 9678 1033
rect 9678 999 9716 1033
rect 9716 999 9750 1033
rect 9750 999 9788 1033
rect 9788 999 9822 1033
rect 9822 999 9855 1033
rect 9611 937 9855 999
rect 9611 903 9644 937
rect 9644 903 9678 937
rect 9678 903 9716 937
rect 9716 903 9750 937
rect 9750 903 9788 937
rect 9788 903 9822 937
rect 9822 903 9855 937
rect 9611 841 9855 903
rect 9611 807 9644 841
rect 9644 807 9678 841
rect 9678 807 9716 841
rect 9716 807 9750 841
rect 9750 807 9788 841
rect 9788 807 9822 841
rect 9822 807 9855 841
rect 9611 745 9855 807
rect 9611 711 9644 745
rect 9644 711 9678 745
rect 9678 711 9716 745
rect 9716 711 9750 745
rect 9750 711 9788 745
rect 9788 711 9822 745
rect 9822 711 9855 745
rect 9611 649 9855 711
rect 9611 615 9644 649
rect 9644 615 9678 649
rect 9678 615 9716 649
rect 9716 615 9750 649
rect 9750 615 9788 649
rect 9788 615 9822 649
rect 9822 615 9855 649
rect 9611 351 9855 615
rect 10023 3337 10267 3382
rect 10023 3303 10056 3337
rect 10056 3303 10090 3337
rect 10090 3303 10128 3337
rect 10128 3303 10162 3337
rect 10162 3303 10200 3337
rect 10200 3303 10234 3337
rect 10234 3303 10267 3337
rect 10023 3241 10267 3303
rect 10023 3207 10056 3241
rect 10056 3207 10090 3241
rect 10090 3207 10128 3241
rect 10128 3207 10162 3241
rect 10162 3207 10200 3241
rect 10200 3207 10234 3241
rect 10234 3207 10267 3241
rect 10023 3145 10267 3207
rect 10023 3111 10056 3145
rect 10056 3111 10090 3145
rect 10090 3111 10128 3145
rect 10128 3111 10162 3145
rect 10162 3111 10200 3145
rect 10200 3111 10234 3145
rect 10234 3111 10267 3145
rect 10023 3049 10267 3111
rect 10023 3015 10056 3049
rect 10056 3015 10090 3049
rect 10090 3015 10128 3049
rect 10128 3015 10162 3049
rect 10162 3015 10200 3049
rect 10200 3015 10234 3049
rect 10234 3015 10267 3049
rect 10023 2953 10267 3015
rect 10023 2919 10056 2953
rect 10056 2919 10090 2953
rect 10090 2919 10128 2953
rect 10128 2919 10162 2953
rect 10162 2919 10200 2953
rect 10200 2919 10234 2953
rect 10234 2919 10267 2953
rect 10023 2857 10267 2919
rect 10023 2823 10056 2857
rect 10056 2823 10090 2857
rect 10090 2823 10128 2857
rect 10128 2823 10162 2857
rect 10162 2823 10200 2857
rect 10200 2823 10234 2857
rect 10234 2823 10267 2857
rect 10023 2761 10267 2823
rect 10023 2727 10056 2761
rect 10056 2727 10090 2761
rect 10090 2727 10128 2761
rect 10128 2727 10162 2761
rect 10162 2727 10200 2761
rect 10200 2727 10234 2761
rect 10234 2727 10267 2761
rect 10023 2665 10267 2727
rect 10023 2631 10056 2665
rect 10056 2631 10090 2665
rect 10090 2631 10128 2665
rect 10128 2631 10162 2665
rect 10162 2631 10200 2665
rect 10200 2631 10234 2665
rect 10234 2631 10267 2665
rect 10023 2569 10267 2631
rect 10023 2535 10056 2569
rect 10056 2535 10090 2569
rect 10090 2535 10128 2569
rect 10128 2535 10162 2569
rect 10162 2535 10200 2569
rect 10200 2535 10234 2569
rect 10234 2535 10267 2569
rect 10023 2473 10267 2535
rect 10023 2439 10056 2473
rect 10056 2439 10090 2473
rect 10090 2439 10128 2473
rect 10128 2439 10162 2473
rect 10162 2439 10200 2473
rect 10200 2439 10234 2473
rect 10234 2439 10267 2473
rect 10023 2377 10267 2439
rect 10023 2343 10056 2377
rect 10056 2343 10090 2377
rect 10090 2343 10128 2377
rect 10128 2343 10162 2377
rect 10162 2343 10200 2377
rect 10200 2343 10234 2377
rect 10234 2343 10267 2377
rect 10023 2281 10267 2343
rect 10023 2247 10056 2281
rect 10056 2247 10090 2281
rect 10090 2247 10128 2281
rect 10128 2247 10162 2281
rect 10162 2247 10200 2281
rect 10200 2247 10234 2281
rect 10234 2247 10267 2281
rect 10023 2185 10267 2247
rect 10023 2151 10056 2185
rect 10056 2151 10090 2185
rect 10090 2151 10128 2185
rect 10128 2151 10162 2185
rect 10162 2151 10200 2185
rect 10200 2151 10234 2185
rect 10234 2151 10267 2185
rect 10023 2089 10267 2151
rect 10023 2055 10056 2089
rect 10056 2055 10090 2089
rect 10090 2055 10128 2089
rect 10128 2055 10162 2089
rect 10162 2055 10200 2089
rect 10200 2055 10234 2089
rect 10234 2055 10267 2089
rect 10023 2050 10267 2055
rect 10435 1863 10468 1875
rect 10468 1863 10502 1875
rect 10502 1863 10540 1875
rect 10540 1863 10574 1875
rect 10574 1863 10612 1875
rect 10612 1863 10646 1875
rect 10646 1863 10679 1875
rect 10435 1801 10679 1863
rect 10435 1767 10468 1801
rect 10468 1767 10502 1801
rect 10502 1767 10540 1801
rect 10540 1767 10574 1801
rect 10574 1767 10612 1801
rect 10612 1767 10646 1801
rect 10646 1767 10679 1801
rect 10435 1705 10679 1767
rect 10435 1671 10468 1705
rect 10468 1671 10502 1705
rect 10502 1671 10540 1705
rect 10540 1671 10574 1705
rect 10574 1671 10612 1705
rect 10612 1671 10646 1705
rect 10646 1671 10679 1705
rect 10435 1609 10679 1671
rect 10435 1575 10468 1609
rect 10468 1575 10502 1609
rect 10502 1575 10540 1609
rect 10540 1575 10574 1609
rect 10574 1575 10612 1609
rect 10612 1575 10646 1609
rect 10646 1575 10679 1609
rect 10435 1513 10679 1575
rect 10435 1479 10468 1513
rect 10468 1479 10502 1513
rect 10502 1479 10540 1513
rect 10540 1479 10574 1513
rect 10574 1479 10612 1513
rect 10612 1479 10646 1513
rect 10646 1479 10679 1513
rect 10435 1417 10679 1479
rect 10435 1383 10468 1417
rect 10468 1383 10502 1417
rect 10502 1383 10540 1417
rect 10540 1383 10574 1417
rect 10574 1383 10612 1417
rect 10612 1383 10646 1417
rect 10646 1383 10679 1417
rect 10435 1321 10679 1383
rect 10435 1287 10468 1321
rect 10468 1287 10502 1321
rect 10502 1287 10540 1321
rect 10540 1287 10574 1321
rect 10574 1287 10612 1321
rect 10612 1287 10646 1321
rect 10646 1287 10679 1321
rect 10435 1225 10679 1287
rect 10435 1191 10468 1225
rect 10468 1191 10502 1225
rect 10502 1191 10540 1225
rect 10540 1191 10574 1225
rect 10574 1191 10612 1225
rect 10612 1191 10646 1225
rect 10646 1191 10679 1225
rect 10435 1129 10679 1191
rect 10435 1095 10468 1129
rect 10468 1095 10502 1129
rect 10502 1095 10540 1129
rect 10540 1095 10574 1129
rect 10574 1095 10612 1129
rect 10612 1095 10646 1129
rect 10646 1095 10679 1129
rect 10435 1033 10679 1095
rect 10435 999 10468 1033
rect 10468 999 10502 1033
rect 10502 999 10540 1033
rect 10540 999 10574 1033
rect 10574 999 10612 1033
rect 10612 999 10646 1033
rect 10646 999 10679 1033
rect 10435 937 10679 999
rect 10435 903 10468 937
rect 10468 903 10502 937
rect 10502 903 10540 937
rect 10540 903 10574 937
rect 10574 903 10612 937
rect 10612 903 10646 937
rect 10646 903 10679 937
rect 10435 841 10679 903
rect 10435 807 10468 841
rect 10468 807 10502 841
rect 10502 807 10540 841
rect 10540 807 10574 841
rect 10574 807 10612 841
rect 10612 807 10646 841
rect 10646 807 10679 841
rect 10435 745 10679 807
rect 10435 711 10468 745
rect 10468 711 10502 745
rect 10502 711 10540 745
rect 10540 711 10574 745
rect 10574 711 10612 745
rect 10612 711 10646 745
rect 10646 711 10679 745
rect 10435 649 10679 711
rect 10435 615 10468 649
rect 10468 615 10502 649
rect 10502 615 10540 649
rect 10540 615 10574 649
rect 10574 615 10612 649
rect 10612 615 10646 649
rect 10646 615 10679 649
rect 10435 351 10679 615
rect 10847 3337 11091 3382
rect 10847 3303 10880 3337
rect 10880 3303 10914 3337
rect 10914 3303 10952 3337
rect 10952 3303 10986 3337
rect 10986 3303 11024 3337
rect 11024 3303 11058 3337
rect 11058 3303 11091 3337
rect 10847 3241 11091 3303
rect 10847 3207 10880 3241
rect 10880 3207 10914 3241
rect 10914 3207 10952 3241
rect 10952 3207 10986 3241
rect 10986 3207 11024 3241
rect 11024 3207 11058 3241
rect 11058 3207 11091 3241
rect 10847 3145 11091 3207
rect 10847 3111 10880 3145
rect 10880 3111 10914 3145
rect 10914 3111 10952 3145
rect 10952 3111 10986 3145
rect 10986 3111 11024 3145
rect 11024 3111 11058 3145
rect 11058 3111 11091 3145
rect 10847 3049 11091 3111
rect 10847 3015 10880 3049
rect 10880 3015 10914 3049
rect 10914 3015 10952 3049
rect 10952 3015 10986 3049
rect 10986 3015 11024 3049
rect 11024 3015 11058 3049
rect 11058 3015 11091 3049
rect 10847 2953 11091 3015
rect 10847 2919 10880 2953
rect 10880 2919 10914 2953
rect 10914 2919 10952 2953
rect 10952 2919 10986 2953
rect 10986 2919 11024 2953
rect 11024 2919 11058 2953
rect 11058 2919 11091 2953
rect 10847 2857 11091 2919
rect 10847 2823 10880 2857
rect 10880 2823 10914 2857
rect 10914 2823 10952 2857
rect 10952 2823 10986 2857
rect 10986 2823 11024 2857
rect 11024 2823 11058 2857
rect 11058 2823 11091 2857
rect 10847 2761 11091 2823
rect 10847 2727 10880 2761
rect 10880 2727 10914 2761
rect 10914 2727 10952 2761
rect 10952 2727 10986 2761
rect 10986 2727 11024 2761
rect 11024 2727 11058 2761
rect 11058 2727 11091 2761
rect 10847 2665 11091 2727
rect 10847 2631 10880 2665
rect 10880 2631 10914 2665
rect 10914 2631 10952 2665
rect 10952 2631 10986 2665
rect 10986 2631 11024 2665
rect 11024 2631 11058 2665
rect 11058 2631 11091 2665
rect 10847 2569 11091 2631
rect 10847 2535 10880 2569
rect 10880 2535 10914 2569
rect 10914 2535 10952 2569
rect 10952 2535 10986 2569
rect 10986 2535 11024 2569
rect 11024 2535 11058 2569
rect 11058 2535 11091 2569
rect 10847 2473 11091 2535
rect 10847 2439 10880 2473
rect 10880 2439 10914 2473
rect 10914 2439 10952 2473
rect 10952 2439 10986 2473
rect 10986 2439 11024 2473
rect 11024 2439 11058 2473
rect 11058 2439 11091 2473
rect 10847 2377 11091 2439
rect 10847 2343 10880 2377
rect 10880 2343 10914 2377
rect 10914 2343 10952 2377
rect 10952 2343 10986 2377
rect 10986 2343 11024 2377
rect 11024 2343 11058 2377
rect 11058 2343 11091 2377
rect 10847 2281 11091 2343
rect 10847 2247 10880 2281
rect 10880 2247 10914 2281
rect 10914 2247 10952 2281
rect 10952 2247 10986 2281
rect 10986 2247 11024 2281
rect 11024 2247 11058 2281
rect 11058 2247 11091 2281
rect 10847 2185 11091 2247
rect 10847 2151 10880 2185
rect 10880 2151 10914 2185
rect 10914 2151 10952 2185
rect 10952 2151 10986 2185
rect 10986 2151 11024 2185
rect 11024 2151 11058 2185
rect 11058 2151 11091 2185
rect 10847 2089 11091 2151
rect 10847 2055 10880 2089
rect 10880 2055 10914 2089
rect 10914 2055 10952 2089
rect 10952 2055 10986 2089
rect 10986 2055 11024 2089
rect 11024 2055 11058 2089
rect 11058 2055 11091 2089
rect 10847 2050 11091 2055
rect 7232 -20 10676 288
<< metal2 >>
rect 7085 3684 10869 3714
rect 7085 3568 7220 3684
rect 10856 3568 10869 3684
rect 7085 3538 10869 3568
rect 7085 3382 11119 3416
rect 7085 2050 7551 3382
rect 7795 2050 8375 3382
rect 8619 2050 9199 3382
rect 9443 2050 10023 3382
rect 10267 2050 10847 3382
rect 11091 2050 11119 3382
rect 7085 2016 11119 2050
rect 7085 1875 11141 1908
rect 7085 351 7963 1875
rect 8207 351 8787 1875
rect 9031 351 9611 1875
rect 9855 351 10435 1875
rect 10679 351 11141 1875
rect 7085 288 11141 351
rect 7085 -20 7232 288
rect 10676 -20 11141 288
rect 7085 -48 11141 -20
<< properties >>
string GDS_END 521198
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 262634
<< end >>
