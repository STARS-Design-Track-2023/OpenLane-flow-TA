* NGSPICE file created from sky130_fd_pr__rf_pnp_05v5_W0p68L0p68.ext - technology: sky130B

.subckt sky130_fd_pr__rf_pnp_05v5_W0p68L0p68 Base Collector Emitter
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0.945
.ends

