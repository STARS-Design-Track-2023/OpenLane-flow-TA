magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -66 377 2850 897
<< pwell >>
rect 2073 287 2780 315
rect 4 221 422 222
rect 1159 221 1417 287
rect 1807 221 2780 287
rect 4 43 2780 221
rect -26 -43 2810 43
<< mvnmos >>
rect 83 112 183 196
rect 239 112 339 196
rect 609 111 709 195
rect 765 111 865 195
rect 921 111 1021 195
rect 1063 111 1163 195
rect 1238 111 1338 261
rect 1413 111 1513 195
rect 1569 111 1669 195
rect 1711 111 1811 195
rect 1886 111 1986 261
rect 2152 139 2252 289
rect 2422 205 2522 289
rect 2601 139 2701 289
<< mvpmos >>
rect 87 488 187 638
rect 243 488 343 638
rect 609 539 709 623
rect 765 539 865 623
rect 921 539 1021 623
rect 1063 539 1163 623
rect 1238 539 1338 739
rect 1394 539 1494 739
rect 1569 539 1669 623
rect 1711 539 1811 623
rect 1886 539 1986 739
rect 2152 443 2252 743
rect 2418 443 2518 593
rect 2597 443 2697 743
<< mvndiff >>
rect 30 171 83 196
rect 30 137 38 171
rect 72 137 83 171
rect 30 112 83 137
rect 183 171 239 196
rect 183 137 194 171
rect 228 137 239 171
rect 183 112 239 137
rect 339 171 396 196
rect 1185 195 1238 261
rect 339 137 350 171
rect 384 137 396 171
rect 339 112 396 137
rect 536 170 609 195
rect 536 136 548 170
rect 582 136 609 170
rect 536 111 609 136
rect 709 172 765 195
rect 709 138 720 172
rect 754 138 765 172
rect 709 111 765 138
rect 865 172 921 195
rect 865 138 876 172
rect 910 138 921 172
rect 865 111 921 138
rect 1021 111 1063 195
rect 1163 177 1238 195
rect 1163 143 1193 177
rect 1227 143 1238 177
rect 1163 111 1238 143
rect 1338 249 1391 261
rect 1338 215 1349 249
rect 1383 215 1391 249
rect 1338 195 1391 215
rect 2099 277 2152 289
rect 1833 249 1886 261
rect 1833 215 1841 249
rect 1875 215 1886 249
rect 1833 195 1886 215
rect 1338 157 1413 195
rect 1338 123 1349 157
rect 1383 123 1413 157
rect 1338 111 1413 123
rect 1513 170 1569 195
rect 1513 136 1524 170
rect 1558 136 1569 170
rect 1513 111 1569 136
rect 1669 111 1711 195
rect 1811 157 1886 195
rect 1811 123 1841 157
rect 1875 123 1886 157
rect 1811 111 1886 123
rect 1986 249 2039 261
rect 1986 215 1997 249
rect 2031 215 2039 249
rect 1986 157 2039 215
rect 1986 123 1997 157
rect 2031 123 2039 157
rect 2099 243 2107 277
rect 2141 243 2152 277
rect 2099 185 2152 243
rect 2099 151 2107 185
rect 2141 151 2152 185
rect 2099 139 2152 151
rect 2252 281 2309 289
rect 2252 247 2263 281
rect 2297 247 2309 281
rect 2252 181 2309 247
rect 2369 264 2422 289
rect 2369 230 2377 264
rect 2411 230 2422 264
rect 2369 205 2422 230
rect 2522 281 2601 289
rect 2522 247 2556 281
rect 2590 247 2601 281
rect 2522 205 2601 247
rect 2252 147 2263 181
rect 2297 147 2309 181
rect 2544 181 2601 205
rect 2252 139 2309 147
rect 2544 147 2556 181
rect 2590 147 2601 181
rect 2544 139 2601 147
rect 2701 277 2754 289
rect 2701 243 2712 277
rect 2746 243 2754 277
rect 2701 185 2754 243
rect 2701 151 2712 185
rect 2746 151 2754 185
rect 2701 139 2754 151
rect 1986 111 2039 123
<< mvpdiff >>
rect 1185 727 1238 739
rect 1185 693 1193 727
rect 1227 693 1238 727
rect 30 630 87 638
rect 30 596 42 630
rect 76 596 87 630
rect 30 530 87 596
rect 30 496 42 530
rect 76 496 87 530
rect 30 488 87 496
rect 187 630 243 638
rect 187 596 198 630
rect 232 596 243 630
rect 187 530 243 596
rect 187 496 198 530
rect 232 496 243 530
rect 187 488 243 496
rect 343 630 400 638
rect 343 596 354 630
rect 388 596 400 630
rect 1185 631 1238 693
rect 1185 623 1193 631
rect 343 530 400 596
rect 552 598 609 623
rect 552 564 564 598
rect 598 564 609 598
rect 552 539 609 564
rect 709 598 765 623
rect 709 564 720 598
rect 754 564 765 598
rect 709 539 765 564
rect 865 598 921 623
rect 865 564 876 598
rect 910 564 921 598
rect 865 539 921 564
rect 1021 539 1063 623
rect 1163 597 1193 623
rect 1227 597 1238 631
rect 1163 539 1238 597
rect 1338 675 1394 739
rect 1338 641 1349 675
rect 1383 641 1394 675
rect 1338 581 1394 641
rect 1338 547 1349 581
rect 1383 547 1394 581
rect 1338 539 1394 547
rect 1494 691 1547 739
rect 1494 657 1505 691
rect 1539 657 1547 691
rect 1494 623 1547 657
rect 1833 727 1886 739
rect 1833 693 1841 727
rect 1875 693 1886 727
rect 1833 656 1886 693
rect 1833 623 1841 656
rect 1494 585 1569 623
rect 1494 551 1505 585
rect 1539 551 1569 585
rect 1494 539 1569 551
rect 1669 539 1711 623
rect 1811 622 1841 623
rect 1875 622 1886 656
rect 1811 585 1886 622
rect 1811 551 1841 585
rect 1875 551 1886 585
rect 1811 539 1886 551
rect 1986 727 2039 739
rect 1986 693 1997 727
rect 2031 693 2039 727
rect 1986 656 2039 693
rect 1986 622 1997 656
rect 2031 622 2039 656
rect 1986 585 2039 622
rect 1986 551 1997 585
rect 2031 551 2039 585
rect 1986 539 2039 551
rect 2099 731 2152 743
rect 2099 697 2107 731
rect 2141 697 2152 731
rect 2099 651 2152 697
rect 2099 617 2107 651
rect 2141 617 2152 651
rect 2099 569 2152 617
rect 343 496 354 530
rect 388 496 400 530
rect 343 488 400 496
rect 2099 535 2107 569
rect 2141 535 2152 569
rect 2099 489 2152 535
rect 2099 455 2107 489
rect 2141 455 2152 489
rect 2099 443 2152 455
rect 2252 731 2305 743
rect 2252 697 2263 731
rect 2297 697 2305 731
rect 2252 651 2305 697
rect 2252 617 2263 651
rect 2297 617 2305 651
rect 2540 735 2597 743
rect 2540 701 2552 735
rect 2586 701 2597 735
rect 2540 652 2597 701
rect 2252 569 2305 617
rect 2540 618 2552 652
rect 2586 618 2597 652
rect 2540 593 2597 618
rect 2252 535 2263 569
rect 2297 535 2305 569
rect 2252 489 2305 535
rect 2252 455 2263 489
rect 2297 455 2305 489
rect 2252 443 2305 455
rect 2365 581 2418 593
rect 2365 547 2373 581
rect 2407 547 2418 581
rect 2365 489 2418 547
rect 2365 455 2373 489
rect 2407 455 2418 489
rect 2365 443 2418 455
rect 2518 568 2597 593
rect 2518 534 2552 568
rect 2586 534 2597 568
rect 2518 485 2597 534
rect 2518 451 2552 485
rect 2586 451 2597 485
rect 2518 443 2597 451
rect 2697 735 2754 743
rect 2697 701 2708 735
rect 2742 701 2754 735
rect 2697 652 2754 701
rect 2697 618 2708 652
rect 2742 618 2754 652
rect 2697 568 2754 618
rect 2697 534 2708 568
rect 2742 534 2754 568
rect 2697 485 2754 534
rect 2697 451 2708 485
rect 2742 451 2754 485
rect 2697 443 2754 451
<< mvndiffc >>
rect 38 137 72 171
rect 194 137 228 171
rect 350 137 384 171
rect 548 136 582 170
rect 720 138 754 172
rect 876 138 910 172
rect 1193 143 1227 177
rect 1349 215 1383 249
rect 1841 215 1875 249
rect 1349 123 1383 157
rect 1524 136 1558 170
rect 1841 123 1875 157
rect 1997 215 2031 249
rect 1997 123 2031 157
rect 2107 243 2141 277
rect 2107 151 2141 185
rect 2263 247 2297 281
rect 2377 230 2411 264
rect 2556 247 2590 281
rect 2263 147 2297 181
rect 2556 147 2590 181
rect 2712 243 2746 277
rect 2712 151 2746 185
<< mvpdiffc >>
rect 1193 693 1227 727
rect 42 596 76 630
rect 42 496 76 530
rect 198 596 232 630
rect 198 496 232 530
rect 354 596 388 630
rect 564 564 598 598
rect 720 564 754 598
rect 876 564 910 598
rect 1193 597 1227 631
rect 1349 641 1383 675
rect 1349 547 1383 581
rect 1505 657 1539 691
rect 1841 693 1875 727
rect 1505 551 1539 585
rect 1841 622 1875 656
rect 1841 551 1875 585
rect 1997 693 2031 727
rect 1997 622 2031 656
rect 1997 551 2031 585
rect 2107 697 2141 731
rect 2107 617 2141 651
rect 354 496 388 530
rect 2107 535 2141 569
rect 2107 455 2141 489
rect 2263 697 2297 731
rect 2263 617 2297 651
rect 2552 701 2586 735
rect 2552 618 2586 652
rect 2263 535 2297 569
rect 2263 455 2297 489
rect 2373 547 2407 581
rect 2373 455 2407 489
rect 2552 534 2586 568
rect 2552 451 2586 485
rect 2708 701 2742 735
rect 2708 618 2742 652
rect 2708 534 2742 568
rect 2708 451 2742 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2784 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
<< poly >>
rect 1238 739 1338 765
rect 1394 739 1494 765
rect 1886 739 1986 765
rect 2152 743 2252 769
rect 2597 743 2697 769
rect 87 638 187 664
rect 243 638 343 664
rect 609 623 709 649
rect 765 623 865 649
rect 921 623 1021 649
rect 1063 623 1163 649
rect 1569 623 1669 649
rect 1711 623 1811 649
rect 87 462 187 488
rect 83 428 187 462
rect 83 394 128 428
rect 162 394 187 428
rect 83 360 187 394
rect 243 378 343 488
rect 609 438 709 539
rect 83 326 128 360
rect 162 326 187 360
rect 83 306 187 326
rect 239 358 343 378
rect 239 324 259 358
rect 293 324 343 358
rect 83 196 183 306
rect 239 290 343 324
rect 239 256 259 290
rect 293 256 343 290
rect 239 222 343 256
rect 600 418 709 438
rect 600 384 620 418
rect 654 384 709 418
rect 765 437 865 539
rect 921 491 1021 539
rect 921 479 967 491
rect 951 457 967 479
rect 1001 457 1021 491
rect 951 441 1021 457
rect 1063 488 1163 539
rect 1063 454 1103 488
rect 1137 454 1163 488
rect 765 399 909 437
rect 600 350 709 384
rect 600 316 620 350
rect 654 316 709 350
rect 239 196 339 222
rect 600 221 709 316
rect 609 195 709 221
rect 751 341 826 357
rect 751 307 776 341
rect 810 307 826 341
rect 868 344 1021 399
rect 868 329 946 344
rect 751 287 826 307
rect 921 310 946 329
rect 980 310 1021 344
rect 751 273 865 287
rect 751 239 776 273
rect 810 239 865 273
rect 751 217 865 239
rect 765 195 865 217
rect 921 276 1021 310
rect 921 242 946 276
rect 980 242 1021 276
rect 921 195 1021 242
rect 1063 195 1163 454
rect 1238 421 1338 539
rect 1394 491 1494 539
rect 1569 513 1669 539
rect 1394 457 1435 491
rect 1469 457 1494 491
rect 1394 437 1494 457
rect 1238 387 1258 421
rect 1292 387 1338 421
rect 1563 395 1669 513
rect 1711 436 1811 539
rect 1886 513 1986 539
rect 1875 486 1986 513
rect 1875 452 1895 486
rect 1929 452 1986 486
rect 1711 416 1825 436
rect 1238 353 1338 387
rect 1238 319 1258 353
rect 1292 319 1338 353
rect 1238 261 1338 319
rect 1413 357 1663 395
rect 1413 323 1445 357
rect 1479 333 1663 357
rect 1711 382 1771 416
rect 1805 382 1825 416
rect 1711 348 1825 382
rect 1875 418 1986 452
rect 2418 593 2518 619
rect 1875 384 1895 418
rect 1929 384 1986 418
rect 2152 417 2252 443
rect 2418 417 2518 443
rect 2597 417 2697 443
rect 1875 364 1986 384
rect 1479 323 1513 333
rect 1413 289 1513 323
rect 1711 314 1771 348
rect 1805 314 1825 348
rect 1711 294 1825 314
rect 83 86 183 112
rect 239 86 339 112
rect 1413 255 1445 289
rect 1479 255 1513 289
rect 1413 195 1513 255
rect 1563 271 1669 291
rect 1563 237 1605 271
rect 1639 237 1669 271
rect 1563 217 1669 237
rect 1569 195 1669 217
rect 1711 195 1811 294
rect 1886 261 1986 364
rect 2031 379 2522 417
rect 2031 345 2051 379
rect 2085 345 2522 379
rect 2031 315 2522 345
rect 2590 383 2701 417
rect 2590 349 2610 383
rect 2644 349 2701 383
rect 2590 315 2701 349
rect 2152 289 2252 315
rect 2422 289 2522 315
rect 2601 289 2701 315
rect 2422 179 2522 205
rect 2152 113 2252 139
rect 2601 113 2701 139
rect 609 85 709 111
rect 765 85 865 111
rect 921 85 1021 111
rect 1063 85 1163 111
rect 1238 85 1338 111
rect 1413 85 1513 111
rect 1569 85 1669 111
rect 1711 85 1811 111
rect 1886 85 1986 111
<< polycont >>
rect 128 394 162 428
rect 128 326 162 360
rect 259 324 293 358
rect 259 256 293 290
rect 620 384 654 418
rect 967 457 1001 491
rect 1103 454 1137 488
rect 620 316 654 350
rect 776 307 810 341
rect 946 310 980 344
rect 776 239 810 273
rect 946 242 980 276
rect 1435 457 1469 491
rect 1258 387 1292 421
rect 1895 452 1929 486
rect 1258 319 1292 353
rect 1445 323 1479 357
rect 1771 382 1805 416
rect 1895 384 1929 418
rect 1771 314 1805 348
rect 1445 255 1479 289
rect 1605 237 1639 271
rect 2051 345 2085 379
rect 2610 349 2644 383
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2784 831
rect 114 735 232 741
rect 114 701 120 735
rect 154 701 192 735
rect 226 701 232 735
rect 494 735 600 741
rect 22 630 76 646
rect 22 596 42 630
rect 22 530 76 596
rect 22 496 42 530
rect 22 274 76 496
rect 114 630 232 701
rect 114 596 198 630
rect 114 530 232 596
rect 114 496 198 530
rect 114 480 232 496
rect 268 682 458 716
rect 112 428 178 444
rect 112 394 128 428
rect 162 394 178 428
rect 112 360 178 394
rect 268 374 302 682
rect 338 630 388 646
rect 338 596 354 630
rect 338 530 388 596
rect 338 496 354 530
rect 338 480 388 496
rect 112 326 128 360
rect 162 326 178 360
rect 112 310 178 326
rect 243 358 309 374
rect 243 324 259 358
rect 293 324 309 358
rect 243 290 309 324
rect 243 274 259 290
rect 22 256 259 274
rect 293 256 309 290
rect 22 240 309 256
rect 350 273 388 480
rect 424 495 458 682
rect 528 701 566 735
rect 1053 735 1243 743
rect 1053 701 1059 735
rect 1093 701 1131 735
rect 1165 727 1203 735
rect 1165 701 1193 727
rect 1237 701 1243 735
rect 494 598 600 701
rect 494 564 564 598
rect 598 564 600 598
rect 494 531 600 564
rect 636 667 1017 701
rect 636 495 670 667
rect 424 461 670 495
rect 706 598 754 631
rect 706 564 720 598
rect 706 531 754 564
rect 505 418 670 425
rect 505 384 620 418
rect 654 384 670 418
rect 505 350 670 384
rect 505 316 620 350
rect 654 316 670 350
rect 505 309 670 316
rect 22 171 88 240
rect 350 239 668 273
rect 22 137 38 171
rect 72 137 88 171
rect 22 108 88 137
rect 124 171 314 204
rect 124 137 194 171
rect 228 137 314 171
rect 124 113 314 137
rect 124 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 314 113
rect 350 171 384 239
rect 350 104 384 137
rect 420 170 598 203
rect 420 136 548 170
rect 582 136 598 170
rect 420 113 598 136
rect 124 73 314 79
rect 454 79 492 113
rect 526 79 564 113
rect 420 73 598 79
rect 634 87 668 239
rect 706 187 740 531
rect 790 357 824 667
rect 776 341 824 357
rect 810 307 824 341
rect 776 273 824 307
rect 810 239 824 273
rect 776 223 824 239
rect 860 598 910 631
rect 860 564 876 598
rect 860 415 910 564
rect 951 561 1017 667
rect 1053 693 1193 701
rect 1227 693 1243 701
rect 1053 631 1243 693
rect 1053 597 1193 631
rect 1227 597 1243 631
rect 1279 727 1649 761
rect 1279 561 1313 727
rect 951 527 1313 561
rect 1349 675 1383 691
rect 1349 581 1383 641
rect 951 491 1017 527
rect 1349 491 1383 547
rect 951 457 967 491
rect 1001 457 1017 491
rect 951 451 1017 457
rect 1087 488 1383 491
rect 1087 454 1103 488
rect 1137 457 1383 488
rect 1137 454 1153 457
rect 1087 451 1153 454
rect 1242 415 1258 421
rect 860 387 1258 415
rect 1292 387 1308 421
rect 860 381 1308 387
rect 860 203 894 381
rect 1242 353 1308 381
rect 930 344 996 345
rect 930 310 946 344
rect 980 310 996 344
rect 1242 319 1258 353
rect 1292 319 1308 353
rect 930 283 996 310
rect 930 276 1297 283
rect 930 242 946 276
rect 980 249 1297 276
rect 1349 265 1383 457
rect 1419 499 1453 727
rect 1489 657 1505 691
rect 1539 657 1559 691
rect 1489 585 1559 657
rect 1489 551 1505 585
rect 1539 551 1559 585
rect 1489 535 1559 551
rect 1419 491 1485 499
rect 1419 457 1435 491
rect 1469 457 1485 491
rect 1419 441 1485 457
rect 1435 357 1489 373
rect 1435 323 1445 357
rect 1479 323 1489 357
rect 1435 289 1489 323
rect 980 242 996 249
rect 930 239 996 242
rect 704 172 770 187
rect 704 138 720 172
rect 754 138 770 172
rect 704 123 770 138
rect 860 172 926 203
rect 860 138 876 172
rect 910 138 926 172
rect 860 123 926 138
rect 962 87 996 239
rect 634 53 996 87
rect 1037 177 1227 213
rect 1037 143 1193 177
rect 1037 113 1227 143
rect 1037 79 1043 113
rect 1077 79 1115 113
rect 1149 79 1187 113
rect 1221 79 1227 113
rect 1037 73 1227 79
rect 1263 87 1297 249
rect 1333 249 1399 265
rect 1333 215 1349 249
rect 1383 215 1399 249
rect 1333 157 1399 215
rect 1333 123 1349 157
rect 1383 123 1399 157
rect 1435 255 1445 289
rect 1479 255 1489 289
rect 1435 239 1489 255
rect 1435 87 1469 239
rect 1525 203 1559 535
rect 1595 271 1649 727
rect 1701 737 1891 743
rect 1701 703 1707 737
rect 1741 703 1779 737
rect 1813 727 1851 737
rect 1813 703 1841 727
rect 1885 703 1891 737
rect 1701 693 1841 703
rect 1875 693 1891 703
rect 1701 656 1891 693
rect 1701 622 1841 656
rect 1875 622 1891 656
rect 1701 585 1891 622
rect 1701 551 1841 585
rect 1875 551 1891 585
rect 1701 535 1891 551
rect 1981 727 2047 743
rect 1981 693 1997 727
rect 2031 693 2047 727
rect 1981 656 2047 693
rect 1981 622 1997 656
rect 2031 622 2047 656
rect 1981 585 2047 622
rect 1981 551 1997 585
rect 2031 551 2047 585
rect 1595 237 1605 271
rect 1639 237 1649 271
rect 1595 221 1649 237
rect 1685 486 1945 499
rect 1685 465 1895 486
rect 1508 170 1559 203
rect 1508 136 1524 170
rect 1558 137 1559 170
rect 1685 137 1719 465
rect 1879 452 1895 465
rect 1929 452 1945 486
rect 1755 416 1821 429
rect 1755 382 1771 416
rect 1805 382 1821 416
rect 1755 348 1821 382
rect 1879 418 1945 452
rect 1879 384 1895 418
rect 1929 384 1945 418
rect 1879 371 1945 384
rect 1981 395 2047 551
rect 2091 731 2178 747
rect 2091 697 2107 731
rect 2141 697 2178 731
rect 2091 651 2178 697
rect 2091 617 2107 651
rect 2141 617 2178 651
rect 2091 569 2178 617
rect 2091 535 2107 569
rect 2141 535 2178 569
rect 2091 489 2178 535
rect 2091 455 2107 489
rect 2141 455 2178 489
rect 2091 439 2178 455
rect 2214 735 2321 747
rect 2248 731 2286 735
rect 2248 701 2263 731
rect 2320 701 2321 735
rect 2214 697 2263 701
rect 2297 697 2321 701
rect 2214 651 2321 697
rect 2214 617 2263 651
rect 2297 617 2321 651
rect 2214 569 2321 617
rect 2459 735 2649 751
rect 2459 701 2465 735
rect 2499 701 2537 735
rect 2586 701 2609 735
rect 2643 701 2649 735
rect 2459 652 2649 701
rect 2459 618 2552 652
rect 2586 618 2649 652
rect 2214 535 2263 569
rect 2297 535 2321 569
rect 2214 489 2321 535
rect 2214 455 2263 489
rect 2297 455 2321 489
rect 2214 439 2321 455
rect 2357 581 2423 597
rect 2357 547 2373 581
rect 2407 547 2423 581
rect 2357 489 2423 547
rect 2357 455 2373 489
rect 2407 455 2423 489
rect 2357 439 2423 455
rect 1981 379 2101 395
rect 1755 314 1771 348
rect 1805 335 1821 348
rect 1981 345 2051 379
rect 2085 345 2101 379
rect 1981 335 2101 345
rect 1805 329 2101 335
rect 1805 314 2047 329
rect 1755 301 2047 314
rect 1558 136 1719 137
rect 1508 103 1719 136
rect 1755 249 1945 265
rect 1755 215 1841 249
rect 1875 215 1945 249
rect 1755 157 1945 215
rect 1755 123 1841 157
rect 1875 123 1945 157
rect 1755 113 1945 123
rect 1263 53 1469 87
rect 1755 79 1761 113
rect 1795 79 1833 113
rect 1867 79 1905 113
rect 1939 79 1945 113
rect 1981 249 2047 301
rect 2137 293 2178 439
rect 2361 399 2423 439
rect 2459 568 2649 618
rect 2459 534 2552 568
rect 2586 534 2649 568
rect 2459 485 2649 534
rect 2459 451 2552 485
rect 2586 451 2649 485
rect 2459 435 2649 451
rect 2692 735 2762 751
rect 2692 701 2708 735
rect 2742 701 2762 735
rect 2692 652 2762 701
rect 2692 618 2708 652
rect 2742 618 2762 652
rect 2692 568 2762 618
rect 2692 534 2708 568
rect 2742 534 2762 568
rect 2692 485 2762 534
rect 2692 451 2708 485
rect 2742 451 2762 485
rect 2692 435 2762 451
rect 2361 383 2660 399
rect 2361 349 2610 383
rect 2644 349 2660 383
rect 2361 333 2660 349
rect 1981 215 1997 249
rect 2031 215 2047 249
rect 1981 157 2047 215
rect 1981 123 1997 157
rect 2031 123 2047 157
rect 2091 277 2178 293
rect 2091 243 2107 277
rect 2141 243 2178 277
rect 2091 185 2178 243
rect 2091 151 2107 185
rect 2141 151 2178 185
rect 2091 135 2178 151
rect 2214 281 2325 297
rect 2214 247 2263 281
rect 2297 247 2325 281
rect 2214 181 2325 247
rect 2361 264 2427 333
rect 2361 230 2377 264
rect 2411 230 2427 264
rect 2361 201 2427 230
rect 2463 281 2653 297
rect 2463 247 2556 281
rect 2590 247 2653 281
rect 2214 147 2263 181
rect 2297 147 2325 181
rect 1981 107 2047 123
rect 2214 113 2325 147
rect 1755 73 1945 79
rect 2214 79 2216 113
rect 2250 79 2288 113
rect 2322 79 2325 113
rect 2214 73 2325 79
rect 2463 181 2653 247
rect 2463 147 2556 181
rect 2590 147 2653 181
rect 2463 113 2653 147
rect 2696 277 2762 435
rect 2696 243 2712 277
rect 2746 243 2762 277
rect 2696 185 2762 243
rect 2696 151 2712 185
rect 2746 151 2762 185
rect 2696 135 2762 151
rect 2463 79 2469 113
rect 2503 79 2541 113
rect 2575 79 2613 113
rect 2647 79 2653 113
rect 2463 73 2653 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 120 701 154 735
rect 192 701 226 735
rect 494 701 528 735
rect 566 701 600 735
rect 1059 701 1093 735
rect 1131 701 1165 735
rect 1203 727 1237 735
rect 1203 701 1227 727
rect 1227 701 1237 727
rect 130 79 164 113
rect 202 79 236 113
rect 274 79 308 113
rect 420 79 454 113
rect 492 79 526 113
rect 564 79 598 113
rect 1043 79 1077 113
rect 1115 79 1149 113
rect 1187 79 1221 113
rect 1707 703 1741 737
rect 1779 703 1813 737
rect 1851 727 1885 737
rect 1851 703 1875 727
rect 1875 703 1885 727
rect 2214 701 2248 735
rect 2286 731 2320 735
rect 2286 701 2297 731
rect 2297 701 2320 731
rect 2465 701 2499 735
rect 2537 701 2552 735
rect 2552 701 2571 735
rect 2609 701 2643 735
rect 1761 79 1795 113
rect 1833 79 1867 113
rect 1905 79 1939 113
rect 2216 79 2250 113
rect 2288 79 2322 113
rect 2469 79 2503 113
rect 2541 79 2575 113
rect 2613 79 2647 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 831 2784 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2784 831
rect 0 791 2784 797
rect 0 737 2784 763
rect 0 735 1707 737
rect 0 701 120 735
rect 154 701 192 735
rect 226 701 494 735
rect 528 701 566 735
rect 600 701 1059 735
rect 1093 701 1131 735
rect 1165 701 1203 735
rect 1237 703 1707 735
rect 1741 703 1779 737
rect 1813 703 1851 737
rect 1885 735 2784 737
rect 1885 703 2214 735
rect 1237 701 2214 703
rect 2248 701 2286 735
rect 2320 701 2465 735
rect 2499 701 2537 735
rect 2571 701 2609 735
rect 2643 701 2784 735
rect 0 689 2784 701
rect 0 113 2784 125
rect 0 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 420 113
rect 454 79 492 113
rect 526 79 564 113
rect 598 79 1043 113
rect 1077 79 1115 113
rect 1149 79 1187 113
rect 1221 79 1761 113
rect 1795 79 1833 113
rect 1867 79 1905 113
rect 1939 79 2216 113
rect 2250 79 2288 113
rect 2322 79 2469 113
rect 2503 79 2541 113
rect 2575 79 2613 113
rect 2647 79 2784 113
rect 0 51 2784 79
rect 0 17 2784 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -23 2784 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfxbp_1
flabel metal1 s 0 51 2784 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 2784 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 689 2784 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 791 2784 814 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2719 242 2753 276 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2719 316 2753 350 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2719 390 2753 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2719 464 2753 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2719 538 2753 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2719 612 2753 646 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2143 168 2177 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2143 242 2177 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2143 316 2177 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2143 390 2177 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2143 464 2177 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2143 538 2177 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2143 612 2177 646 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2784 814
string GDS_END 889718
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 861306
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
