magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 3 21 735 203
rect 28 -17 62 21
<< locali >>
rect 17 214 87 493
rect 17 51 71 214
rect 304 265 358 414
rect 189 199 256 265
rect 290 199 358 265
rect 396 265 443 414
rect 396 199 454 265
rect 488 199 568 265
rect 670 199 719 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 121 367 202 527
rect 236 459 543 493
rect 236 333 270 459
rect 121 299 270 333
rect 121 199 155 299
rect 477 333 543 459
rect 580 367 627 527
rect 661 333 719 493
rect 477 299 719 333
rect 602 165 636 299
rect 105 17 239 165
rect 273 131 552 165
rect 273 62 332 131
rect 368 17 443 97
rect 486 62 552 131
rect 602 51 719 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 189 199 256 265 6 A1
port 1 nsew signal input
rlabel locali s 290 199 358 265 6 A2
port 2 nsew signal input
rlabel locali s 304 265 358 414 6 A2
port 2 nsew signal input
rlabel locali s 396 199 454 265 6 A3
port 3 nsew signal input
rlabel locali s 396 265 443 414 6 A3
port 3 nsew signal input
rlabel locali s 488 199 568 265 6 B1
port 4 nsew signal input
rlabel locali s 670 199 719 265 6 C1
port 5 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 28 -17 62 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 3 21 735 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 17 51 71 214 6 X
port 10 nsew signal output
rlabel locali s 17 214 87 493 6 X
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 920548
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 912932
<< end >>
