magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< metal4 >>
rect 8 39952 15008 39987
rect 8 39716 249 39952
rect 485 39716 576 39952
rect 812 39716 903 39952
rect 1139 39716 1230 39952
rect 1466 39716 1557 39952
rect 1793 39716 1884 39952
rect 2120 39716 2211 39952
rect 2447 39716 2538 39952
rect 2774 39716 2865 39952
rect 3101 39716 3192 39952
rect 3428 39716 3519 39952
rect 3755 39716 3846 39952
rect 4082 39716 4173 39952
rect 4409 39716 4500 39952
rect 4736 39716 4827 39952
rect 5063 39716 5154 39952
rect 5390 39716 5481 39952
rect 5717 39716 5808 39952
rect 6044 39716 6135 39952
rect 6371 39716 6462 39952
rect 6698 39716 6789 39952
rect 7025 39716 7116 39952
rect 7352 39716 7443 39952
rect 7679 39716 7770 39952
rect 8006 39716 8097 39952
rect 8333 39716 8423 39952
rect 8659 39716 8749 39952
rect 8985 39716 9075 39952
rect 9311 39716 9401 39952
rect 9637 39716 9727 39952
rect 9963 39716 10053 39952
rect 10289 39716 10379 39952
rect 10615 39716 10705 39952
rect 10941 39716 11031 39952
rect 11267 39716 11357 39952
rect 11593 39716 11683 39952
rect 11919 39716 12009 39952
rect 12245 39716 12335 39952
rect 12571 39716 12661 39952
rect 12897 39716 12987 39952
rect 13223 39716 13313 39952
rect 13549 39716 13639 39952
rect 13875 39716 13965 39952
rect 14201 39716 14291 39952
rect 14527 39716 14617 39952
rect 14853 39716 15008 39952
rect 8 39628 15008 39716
rect 8 39392 249 39628
rect 485 39392 576 39628
rect 812 39392 903 39628
rect 1139 39392 1230 39628
rect 1466 39392 1557 39628
rect 1793 39392 1884 39628
rect 2120 39392 2211 39628
rect 2447 39392 2538 39628
rect 2774 39392 2865 39628
rect 3101 39392 3192 39628
rect 3428 39392 3519 39628
rect 3755 39392 3846 39628
rect 4082 39392 4173 39628
rect 4409 39392 4500 39628
rect 4736 39392 4827 39628
rect 5063 39392 5154 39628
rect 5390 39392 5481 39628
rect 5717 39392 5808 39628
rect 6044 39392 6135 39628
rect 6371 39392 6462 39628
rect 6698 39392 6789 39628
rect 7025 39392 7116 39628
rect 7352 39392 7443 39628
rect 7679 39392 7770 39628
rect 8006 39392 8097 39628
rect 8333 39392 8423 39628
rect 8659 39392 8749 39628
rect 8985 39392 9075 39628
rect 9311 39392 9401 39628
rect 9637 39392 9727 39628
rect 9963 39392 10053 39628
rect 10289 39392 10379 39628
rect 10615 39392 10705 39628
rect 10941 39392 11031 39628
rect 11267 39392 11357 39628
rect 11593 39392 11683 39628
rect 11919 39392 12009 39628
rect 12245 39392 12335 39628
rect 12571 39392 12661 39628
rect 12897 39392 12987 39628
rect 13223 39392 13313 39628
rect 13549 39392 13639 39628
rect 13875 39392 13965 39628
rect 14201 39392 14291 39628
rect 14527 39392 14617 39628
rect 14853 39392 15008 39628
rect 8 39304 15008 39392
rect 8 39068 249 39304
rect 485 39068 576 39304
rect 812 39068 903 39304
rect 1139 39068 1230 39304
rect 1466 39068 1557 39304
rect 1793 39068 1884 39304
rect 2120 39068 2211 39304
rect 2447 39068 2538 39304
rect 2774 39068 2865 39304
rect 3101 39068 3192 39304
rect 3428 39068 3519 39304
rect 3755 39068 3846 39304
rect 4082 39068 4173 39304
rect 4409 39068 4500 39304
rect 4736 39068 4827 39304
rect 5063 39068 5154 39304
rect 5390 39068 5481 39304
rect 5717 39068 5808 39304
rect 6044 39068 6135 39304
rect 6371 39068 6462 39304
rect 6698 39068 6789 39304
rect 7025 39068 7116 39304
rect 7352 39068 7443 39304
rect 7679 39068 7770 39304
rect 8006 39068 8097 39304
rect 8333 39068 8423 39304
rect 8659 39068 8749 39304
rect 8985 39068 9075 39304
rect 9311 39068 9401 39304
rect 9637 39068 9727 39304
rect 9963 39068 10053 39304
rect 10289 39068 10379 39304
rect 10615 39068 10705 39304
rect 10941 39068 11031 39304
rect 11267 39068 11357 39304
rect 11593 39068 11683 39304
rect 11919 39068 12009 39304
rect 12245 39068 12335 39304
rect 12571 39068 12661 39304
rect 12897 39068 12987 39304
rect 13223 39068 13313 39304
rect 13549 39068 13639 39304
rect 13875 39068 13965 39304
rect 14201 39068 14291 39304
rect 14527 39068 14617 39304
rect 14853 39068 15008 39304
rect 8 38980 15008 39068
rect 8 38744 249 38980
rect 485 38744 576 38980
rect 812 38744 903 38980
rect 1139 38744 1230 38980
rect 1466 38744 1557 38980
rect 1793 38744 1884 38980
rect 2120 38744 2211 38980
rect 2447 38744 2538 38980
rect 2774 38744 2865 38980
rect 3101 38744 3192 38980
rect 3428 38744 3519 38980
rect 3755 38744 3846 38980
rect 4082 38744 4173 38980
rect 4409 38744 4500 38980
rect 4736 38744 4827 38980
rect 5063 38744 5154 38980
rect 5390 38744 5481 38980
rect 5717 38744 5808 38980
rect 6044 38744 6135 38980
rect 6371 38744 6462 38980
rect 6698 38744 6789 38980
rect 7025 38744 7116 38980
rect 7352 38744 7443 38980
rect 7679 38744 7770 38980
rect 8006 38744 8097 38980
rect 8333 38744 8423 38980
rect 8659 38744 8749 38980
rect 8985 38744 9075 38980
rect 9311 38744 9401 38980
rect 9637 38744 9727 38980
rect 9963 38744 10053 38980
rect 10289 38744 10379 38980
rect 10615 38744 10705 38980
rect 10941 38744 11031 38980
rect 11267 38744 11357 38980
rect 11593 38744 11683 38980
rect 11919 38744 12009 38980
rect 12245 38744 12335 38980
rect 12571 38744 12661 38980
rect 12897 38744 12987 38980
rect 13223 38744 13313 38980
rect 13549 38744 13639 38980
rect 13875 38744 13965 38980
rect 14201 38744 14291 38980
rect 14527 38744 14617 38980
rect 14853 38744 15008 38980
rect 8 38656 15008 38744
rect 8 38420 249 38656
rect 485 38420 576 38656
rect 812 38420 903 38656
rect 1139 38420 1230 38656
rect 1466 38420 1557 38656
rect 1793 38420 1884 38656
rect 2120 38420 2211 38656
rect 2447 38420 2538 38656
rect 2774 38420 2865 38656
rect 3101 38420 3192 38656
rect 3428 38420 3519 38656
rect 3755 38420 3846 38656
rect 4082 38420 4173 38656
rect 4409 38420 4500 38656
rect 4736 38420 4827 38656
rect 5063 38420 5154 38656
rect 5390 38420 5481 38656
rect 5717 38420 5808 38656
rect 6044 38420 6135 38656
rect 6371 38420 6462 38656
rect 6698 38420 6789 38656
rect 7025 38420 7116 38656
rect 7352 38420 7443 38656
rect 7679 38420 7770 38656
rect 8006 38420 8097 38656
rect 8333 38420 8423 38656
rect 8659 38420 8749 38656
rect 8985 38420 9075 38656
rect 9311 38420 9401 38656
rect 9637 38420 9727 38656
rect 9963 38420 10053 38656
rect 10289 38420 10379 38656
rect 10615 38420 10705 38656
rect 10941 38420 11031 38656
rect 11267 38420 11357 38656
rect 11593 38420 11683 38656
rect 11919 38420 12009 38656
rect 12245 38420 12335 38656
rect 12571 38420 12661 38656
rect 12897 38420 12987 38656
rect 13223 38420 13313 38656
rect 13549 38420 13639 38656
rect 13875 38420 13965 38656
rect 14201 38420 14291 38656
rect 14527 38420 14617 38656
rect 14853 38420 15008 38656
rect 8 38332 15008 38420
rect 8 38096 249 38332
rect 485 38096 576 38332
rect 812 38096 903 38332
rect 1139 38096 1230 38332
rect 1466 38096 1557 38332
rect 1793 38096 1884 38332
rect 2120 38096 2211 38332
rect 2447 38096 2538 38332
rect 2774 38096 2865 38332
rect 3101 38096 3192 38332
rect 3428 38096 3519 38332
rect 3755 38096 3846 38332
rect 4082 38096 4173 38332
rect 4409 38096 4500 38332
rect 4736 38096 4827 38332
rect 5063 38096 5154 38332
rect 5390 38096 5481 38332
rect 5717 38096 5808 38332
rect 6044 38096 6135 38332
rect 6371 38096 6462 38332
rect 6698 38096 6789 38332
rect 7025 38096 7116 38332
rect 7352 38096 7443 38332
rect 7679 38096 7770 38332
rect 8006 38096 8097 38332
rect 8333 38096 8423 38332
rect 8659 38096 8749 38332
rect 8985 38096 9075 38332
rect 9311 38096 9401 38332
rect 9637 38096 9727 38332
rect 9963 38096 10053 38332
rect 10289 38096 10379 38332
rect 10615 38096 10705 38332
rect 10941 38096 11031 38332
rect 11267 38096 11357 38332
rect 11593 38096 11683 38332
rect 11919 38096 12009 38332
rect 12245 38096 12335 38332
rect 12571 38096 12661 38332
rect 12897 38096 12987 38332
rect 13223 38096 13313 38332
rect 13549 38096 13639 38332
rect 13875 38096 13965 38332
rect 14201 38096 14291 38332
rect 14527 38096 14617 38332
rect 14853 38096 15008 38332
rect 8 38008 15008 38096
rect 8 37772 249 38008
rect 485 37772 576 38008
rect 812 37772 903 38008
rect 1139 37772 1230 38008
rect 1466 37772 1557 38008
rect 1793 37772 1884 38008
rect 2120 37772 2211 38008
rect 2447 37772 2538 38008
rect 2774 37772 2865 38008
rect 3101 37772 3192 38008
rect 3428 37772 3519 38008
rect 3755 37772 3846 38008
rect 4082 37772 4173 38008
rect 4409 37772 4500 38008
rect 4736 37772 4827 38008
rect 5063 37772 5154 38008
rect 5390 37772 5481 38008
rect 5717 37772 5808 38008
rect 6044 37772 6135 38008
rect 6371 37772 6462 38008
rect 6698 37772 6789 38008
rect 7025 37772 7116 38008
rect 7352 37772 7443 38008
rect 7679 37772 7770 38008
rect 8006 37772 8097 38008
rect 8333 37772 8423 38008
rect 8659 37772 8749 38008
rect 8985 37772 9075 38008
rect 9311 37772 9401 38008
rect 9637 37772 9727 38008
rect 9963 37772 10053 38008
rect 10289 37772 10379 38008
rect 10615 37772 10705 38008
rect 10941 37772 11031 38008
rect 11267 37772 11357 38008
rect 11593 37772 11683 38008
rect 11919 37772 12009 38008
rect 12245 37772 12335 38008
rect 12571 37772 12661 38008
rect 12897 37772 12987 38008
rect 13223 37772 13313 38008
rect 13549 37772 13639 38008
rect 13875 37772 13965 38008
rect 14201 37772 14291 38008
rect 14527 37772 14617 38008
rect 14853 37772 15008 38008
rect 8 37684 15008 37772
rect 8 37448 249 37684
rect 485 37448 576 37684
rect 812 37448 903 37684
rect 1139 37448 1230 37684
rect 1466 37448 1557 37684
rect 1793 37448 1884 37684
rect 2120 37448 2211 37684
rect 2447 37448 2538 37684
rect 2774 37448 2865 37684
rect 3101 37448 3192 37684
rect 3428 37448 3519 37684
rect 3755 37448 3846 37684
rect 4082 37448 4173 37684
rect 4409 37448 4500 37684
rect 4736 37448 4827 37684
rect 5063 37448 5154 37684
rect 5390 37448 5481 37684
rect 5717 37448 5808 37684
rect 6044 37448 6135 37684
rect 6371 37448 6462 37684
rect 6698 37448 6789 37684
rect 7025 37448 7116 37684
rect 7352 37448 7443 37684
rect 7679 37448 7770 37684
rect 8006 37448 8097 37684
rect 8333 37448 8423 37684
rect 8659 37448 8749 37684
rect 8985 37448 9075 37684
rect 9311 37448 9401 37684
rect 9637 37448 9727 37684
rect 9963 37448 10053 37684
rect 10289 37448 10379 37684
rect 10615 37448 10705 37684
rect 10941 37448 11031 37684
rect 11267 37448 11357 37684
rect 11593 37448 11683 37684
rect 11919 37448 12009 37684
rect 12245 37448 12335 37684
rect 12571 37448 12661 37684
rect 12897 37448 12987 37684
rect 13223 37448 13313 37684
rect 13549 37448 13639 37684
rect 13875 37448 13965 37684
rect 14201 37448 14291 37684
rect 14527 37448 14617 37684
rect 14853 37448 15008 37684
rect 8 37360 15008 37448
rect 8 37124 249 37360
rect 485 37124 576 37360
rect 812 37124 903 37360
rect 1139 37124 1230 37360
rect 1466 37124 1557 37360
rect 1793 37124 1884 37360
rect 2120 37124 2211 37360
rect 2447 37124 2538 37360
rect 2774 37124 2865 37360
rect 3101 37124 3192 37360
rect 3428 37124 3519 37360
rect 3755 37124 3846 37360
rect 4082 37124 4173 37360
rect 4409 37124 4500 37360
rect 4736 37124 4827 37360
rect 5063 37124 5154 37360
rect 5390 37124 5481 37360
rect 5717 37124 5808 37360
rect 6044 37124 6135 37360
rect 6371 37124 6462 37360
rect 6698 37124 6789 37360
rect 7025 37124 7116 37360
rect 7352 37124 7443 37360
rect 7679 37124 7770 37360
rect 8006 37124 8097 37360
rect 8333 37124 8423 37360
rect 8659 37124 8749 37360
rect 8985 37124 9075 37360
rect 9311 37124 9401 37360
rect 9637 37124 9727 37360
rect 9963 37124 10053 37360
rect 10289 37124 10379 37360
rect 10615 37124 10705 37360
rect 10941 37124 11031 37360
rect 11267 37124 11357 37360
rect 11593 37124 11683 37360
rect 11919 37124 12009 37360
rect 12245 37124 12335 37360
rect 12571 37124 12661 37360
rect 12897 37124 12987 37360
rect 13223 37124 13313 37360
rect 13549 37124 13639 37360
rect 13875 37124 13965 37360
rect 14201 37124 14291 37360
rect 14527 37124 14617 37360
rect 14853 37124 15008 37360
rect 8 37036 15008 37124
rect 8 36800 249 37036
rect 485 36800 576 37036
rect 812 36800 903 37036
rect 1139 36800 1230 37036
rect 1466 36800 1557 37036
rect 1793 36800 1884 37036
rect 2120 36800 2211 37036
rect 2447 36800 2538 37036
rect 2774 36800 2865 37036
rect 3101 36800 3192 37036
rect 3428 36800 3519 37036
rect 3755 36800 3846 37036
rect 4082 36800 4173 37036
rect 4409 36800 4500 37036
rect 4736 36800 4827 37036
rect 5063 36800 5154 37036
rect 5390 36800 5481 37036
rect 5717 36800 5808 37036
rect 6044 36800 6135 37036
rect 6371 36800 6462 37036
rect 6698 36800 6789 37036
rect 7025 36800 7116 37036
rect 7352 36800 7443 37036
rect 7679 36800 7770 37036
rect 8006 36800 8097 37036
rect 8333 36800 8423 37036
rect 8659 36800 8749 37036
rect 8985 36800 9075 37036
rect 9311 36800 9401 37036
rect 9637 36800 9727 37036
rect 9963 36800 10053 37036
rect 10289 36800 10379 37036
rect 10615 36800 10705 37036
rect 10941 36800 11031 37036
rect 11267 36800 11357 37036
rect 11593 36800 11683 37036
rect 11919 36800 12009 37036
rect 12245 36800 12335 37036
rect 12571 36800 12661 37036
rect 12897 36800 12987 37036
rect 13223 36800 13313 37036
rect 13549 36800 13639 37036
rect 13875 36800 13965 37036
rect 14201 36800 14291 37036
rect 14527 36800 14617 37036
rect 14853 36800 15008 37036
rect 8 36712 15008 36800
rect 8 36476 249 36712
rect 485 36476 576 36712
rect 812 36476 903 36712
rect 1139 36476 1230 36712
rect 1466 36476 1557 36712
rect 1793 36476 1884 36712
rect 2120 36476 2211 36712
rect 2447 36476 2538 36712
rect 2774 36476 2865 36712
rect 3101 36476 3192 36712
rect 3428 36476 3519 36712
rect 3755 36476 3846 36712
rect 4082 36476 4173 36712
rect 4409 36476 4500 36712
rect 4736 36476 4827 36712
rect 5063 36476 5154 36712
rect 5390 36476 5481 36712
rect 5717 36476 5808 36712
rect 6044 36476 6135 36712
rect 6371 36476 6462 36712
rect 6698 36476 6789 36712
rect 7025 36476 7116 36712
rect 7352 36476 7443 36712
rect 7679 36476 7770 36712
rect 8006 36476 8097 36712
rect 8333 36476 8423 36712
rect 8659 36476 8749 36712
rect 8985 36476 9075 36712
rect 9311 36476 9401 36712
rect 9637 36476 9727 36712
rect 9963 36476 10053 36712
rect 10289 36476 10379 36712
rect 10615 36476 10705 36712
rect 10941 36476 11031 36712
rect 11267 36476 11357 36712
rect 11593 36476 11683 36712
rect 11919 36476 12009 36712
rect 12245 36476 12335 36712
rect 12571 36476 12661 36712
rect 12897 36476 12987 36712
rect 13223 36476 13313 36712
rect 13549 36476 13639 36712
rect 13875 36476 13965 36712
rect 14201 36476 14291 36712
rect 14527 36476 14617 36712
rect 14853 36476 15008 36712
rect 8 36388 15008 36476
rect 8 36152 249 36388
rect 485 36152 576 36388
rect 812 36152 903 36388
rect 1139 36152 1230 36388
rect 1466 36152 1557 36388
rect 1793 36152 1884 36388
rect 2120 36152 2211 36388
rect 2447 36152 2538 36388
rect 2774 36152 2865 36388
rect 3101 36152 3192 36388
rect 3428 36152 3519 36388
rect 3755 36152 3846 36388
rect 4082 36152 4173 36388
rect 4409 36152 4500 36388
rect 4736 36152 4827 36388
rect 5063 36152 5154 36388
rect 5390 36152 5481 36388
rect 5717 36152 5808 36388
rect 6044 36152 6135 36388
rect 6371 36152 6462 36388
rect 6698 36152 6789 36388
rect 7025 36152 7116 36388
rect 7352 36152 7443 36388
rect 7679 36152 7770 36388
rect 8006 36152 8097 36388
rect 8333 36152 8423 36388
rect 8659 36152 8749 36388
rect 8985 36152 9075 36388
rect 9311 36152 9401 36388
rect 9637 36152 9727 36388
rect 9963 36152 10053 36388
rect 10289 36152 10379 36388
rect 10615 36152 10705 36388
rect 10941 36152 11031 36388
rect 11267 36152 11357 36388
rect 11593 36152 11683 36388
rect 11919 36152 12009 36388
rect 12245 36152 12335 36388
rect 12571 36152 12661 36388
rect 12897 36152 12987 36388
rect 13223 36152 13313 36388
rect 13549 36152 13639 36388
rect 13875 36152 13965 36388
rect 14201 36152 14291 36388
rect 14527 36152 14617 36388
rect 14853 36152 15008 36388
rect 8 36064 15008 36152
rect 8 35828 249 36064
rect 485 35828 576 36064
rect 812 35828 903 36064
rect 1139 35828 1230 36064
rect 1466 35828 1557 36064
rect 1793 35828 1884 36064
rect 2120 35828 2211 36064
rect 2447 35828 2538 36064
rect 2774 35828 2865 36064
rect 3101 35828 3192 36064
rect 3428 35828 3519 36064
rect 3755 35828 3846 36064
rect 4082 35828 4173 36064
rect 4409 35828 4500 36064
rect 4736 35828 4827 36064
rect 5063 35828 5154 36064
rect 5390 35828 5481 36064
rect 5717 35828 5808 36064
rect 6044 35828 6135 36064
rect 6371 35828 6462 36064
rect 6698 35828 6789 36064
rect 7025 35828 7116 36064
rect 7352 35828 7443 36064
rect 7679 35828 7770 36064
rect 8006 35828 8097 36064
rect 8333 35828 8423 36064
rect 8659 35828 8749 36064
rect 8985 35828 9075 36064
rect 9311 35828 9401 36064
rect 9637 35828 9727 36064
rect 9963 35828 10053 36064
rect 10289 35828 10379 36064
rect 10615 35828 10705 36064
rect 10941 35828 11031 36064
rect 11267 35828 11357 36064
rect 11593 35828 11683 36064
rect 11919 35828 12009 36064
rect 12245 35828 12335 36064
rect 12571 35828 12661 36064
rect 12897 35828 12987 36064
rect 13223 35828 13313 36064
rect 13549 35828 13639 36064
rect 13875 35828 13965 36064
rect 14201 35828 14291 36064
rect 14527 35828 14617 36064
rect 14853 35828 15008 36064
rect 8 35740 15008 35828
rect 8 35504 249 35740
rect 485 35504 576 35740
rect 812 35504 903 35740
rect 1139 35504 1230 35740
rect 1466 35504 1557 35740
rect 1793 35504 1884 35740
rect 2120 35504 2211 35740
rect 2447 35504 2538 35740
rect 2774 35504 2865 35740
rect 3101 35504 3192 35740
rect 3428 35504 3519 35740
rect 3755 35504 3846 35740
rect 4082 35504 4173 35740
rect 4409 35504 4500 35740
rect 4736 35504 4827 35740
rect 5063 35504 5154 35740
rect 5390 35504 5481 35740
rect 5717 35504 5808 35740
rect 6044 35504 6135 35740
rect 6371 35504 6462 35740
rect 6698 35504 6789 35740
rect 7025 35504 7116 35740
rect 7352 35504 7443 35740
rect 7679 35504 7770 35740
rect 8006 35504 8097 35740
rect 8333 35504 8423 35740
rect 8659 35504 8749 35740
rect 8985 35504 9075 35740
rect 9311 35504 9401 35740
rect 9637 35504 9727 35740
rect 9963 35504 10053 35740
rect 10289 35504 10379 35740
rect 10615 35504 10705 35740
rect 10941 35504 11031 35740
rect 11267 35504 11357 35740
rect 11593 35504 11683 35740
rect 11919 35504 12009 35740
rect 12245 35504 12335 35740
rect 12571 35504 12661 35740
rect 12897 35504 12987 35740
rect 13223 35504 13313 35740
rect 13549 35504 13639 35740
rect 13875 35504 13965 35740
rect 14201 35504 14291 35740
rect 14527 35504 14617 35740
rect 14853 35504 15008 35740
rect 8 35416 15008 35504
rect 8 35180 249 35416
rect 485 35180 576 35416
rect 812 35180 903 35416
rect 1139 35180 1230 35416
rect 1466 35180 1557 35416
rect 1793 35180 1884 35416
rect 2120 35180 2211 35416
rect 2447 35180 2538 35416
rect 2774 35180 2865 35416
rect 3101 35180 3192 35416
rect 3428 35180 3519 35416
rect 3755 35180 3846 35416
rect 4082 35180 4173 35416
rect 4409 35180 4500 35416
rect 4736 35180 4827 35416
rect 5063 35180 5154 35416
rect 5390 35180 5481 35416
rect 5717 35180 5808 35416
rect 6044 35180 6135 35416
rect 6371 35180 6462 35416
rect 6698 35180 6789 35416
rect 7025 35180 7116 35416
rect 7352 35180 7443 35416
rect 7679 35180 7770 35416
rect 8006 35180 8097 35416
rect 8333 35180 8423 35416
rect 8659 35180 8749 35416
rect 8985 35180 9075 35416
rect 9311 35180 9401 35416
rect 9637 35180 9727 35416
rect 9963 35180 10053 35416
rect 10289 35180 10379 35416
rect 10615 35180 10705 35416
rect 10941 35180 11031 35416
rect 11267 35180 11357 35416
rect 11593 35180 11683 35416
rect 11919 35180 12009 35416
rect 12245 35180 12335 35416
rect 12571 35180 12661 35416
rect 12897 35180 12987 35416
rect 13223 35180 13313 35416
rect 13549 35180 13639 35416
rect 13875 35180 13965 35416
rect 14201 35180 14291 35416
rect 14527 35180 14617 35416
rect 14853 35180 15008 35416
rect 8 35144 15008 35180
rect 8 18959 5630 18987
rect 8 18723 151 18959
rect 387 18723 473 18959
rect 709 18723 795 18959
rect 1031 18723 1117 18959
rect 1353 18723 1439 18959
rect 1675 18723 1761 18959
rect 1997 18723 2083 18959
rect 2319 18723 2405 18959
rect 2641 18723 2727 18959
rect 2963 18723 3049 18959
rect 3285 18723 3371 18959
rect 3607 18723 3693 18959
rect 3929 18723 4015 18959
rect 4251 18723 4337 18959
rect 4573 18723 4659 18959
rect 4895 18723 4981 18959
rect 5217 18723 5303 18959
rect 5539 18787 5630 18959
tri 5630 18787 5830 18987 sw
rect 5539 18723 5830 18787
rect 8 18623 5830 18723
rect 8 18387 151 18623
rect 387 18387 473 18623
rect 709 18387 795 18623
rect 1031 18387 1117 18623
rect 1353 18387 1439 18623
rect 1675 18387 1761 18623
rect 1997 18387 2083 18623
rect 2319 18387 2405 18623
rect 2641 18387 2727 18623
rect 2963 18387 3049 18623
rect 3285 18387 3371 18623
rect 3607 18387 3693 18623
rect 3929 18387 4015 18623
rect 4251 18387 4337 18623
rect 4573 18387 4659 18623
rect 4895 18387 4981 18623
rect 5217 18387 5303 18623
rect 5539 18387 5830 18623
rect 8 18287 5830 18387
rect 8 18051 151 18287
rect 387 18051 473 18287
rect 709 18051 795 18287
rect 1031 18051 1117 18287
rect 1353 18051 1439 18287
rect 1675 18051 1761 18287
rect 1997 18051 2083 18287
rect 2319 18051 2405 18287
rect 2641 18051 2727 18287
rect 2963 18051 3049 18287
rect 3285 18051 3371 18287
rect 3607 18051 3693 18287
rect 3929 18051 4015 18287
rect 4251 18051 4337 18287
rect 4573 18051 4659 18287
rect 4895 18051 4981 18287
rect 5217 18051 5303 18287
rect 5539 18051 5830 18287
rect 8 17951 5830 18051
rect 8 17715 151 17951
rect 387 17715 473 17951
rect 709 17715 795 17951
rect 1031 17715 1117 17951
rect 1353 17715 1439 17951
rect 1675 17715 1761 17951
rect 1997 17715 2083 17951
rect 2319 17715 2405 17951
rect 2641 17715 2727 17951
rect 2963 17715 3049 17951
rect 3285 17715 3371 17951
rect 3607 17715 3693 17951
rect 3929 17715 4015 17951
rect 4251 17715 4337 17951
rect 4573 17715 4659 17951
rect 4895 17715 4981 17951
rect 5217 17715 5303 17951
rect 5539 17715 5830 17951
rect 8 17615 5830 17715
rect 8 17379 151 17615
rect 387 17379 473 17615
rect 709 17379 795 17615
rect 1031 17379 1117 17615
rect 1353 17379 1439 17615
rect 1675 17379 1761 17615
rect 1997 17379 2083 17615
rect 2319 17379 2405 17615
rect 2641 17379 2727 17615
rect 2963 17379 3049 17615
rect 3285 17379 3371 17615
rect 3607 17379 3693 17615
rect 3929 17379 4015 17615
rect 4251 17379 4337 17615
rect 4573 17379 4659 17615
rect 4895 17379 4981 17615
rect 5217 17379 5303 17615
rect 5539 17379 5830 17615
rect 8 17279 5830 17379
rect 8 17043 151 17279
rect 387 17043 473 17279
rect 709 17043 795 17279
rect 1031 17043 1117 17279
rect 1353 17043 1439 17279
rect 1675 17043 1761 17279
rect 1997 17043 2083 17279
rect 2319 17043 2405 17279
rect 2641 17043 2727 17279
rect 2963 17043 3049 17279
rect 3285 17043 3371 17279
rect 3607 17043 3693 17279
rect 3929 17043 4015 17279
rect 4251 17043 4337 17279
rect 4573 17043 4659 17279
rect 4895 17043 4981 17279
rect 5217 17043 5303 17279
rect 5539 17043 5830 17279
rect 8 16943 5830 17043
rect 8 16707 151 16943
rect 387 16707 473 16943
rect 709 16707 795 16943
rect 1031 16707 1117 16943
rect 1353 16707 1439 16943
rect 1675 16707 1761 16943
rect 1997 16707 2083 16943
rect 2319 16707 2405 16943
rect 2641 16707 2727 16943
rect 2963 16707 3049 16943
rect 3285 16707 3371 16943
rect 3607 16707 3693 16943
rect 3929 16707 4015 16943
rect 4251 16707 4337 16943
rect 4573 16707 4659 16943
rect 4895 16707 4981 16943
rect 5217 16707 5303 16943
rect 5539 16707 5830 16943
rect 8 16607 5830 16707
rect 8 16371 151 16607
rect 387 16371 473 16607
rect 709 16371 795 16607
rect 1031 16371 1117 16607
rect 1353 16371 1439 16607
rect 1675 16371 1761 16607
rect 1997 16371 2083 16607
rect 2319 16371 2405 16607
rect 2641 16371 2727 16607
rect 2963 16371 3049 16607
rect 3285 16371 3371 16607
rect 3607 16371 3693 16607
rect 3929 16371 4015 16607
rect 4251 16371 4337 16607
rect 4573 16371 4659 16607
rect 4895 16371 4981 16607
rect 5217 16371 5303 16607
rect 5539 16371 5830 16607
rect 8 16271 5830 16371
rect 8 16035 151 16271
rect 387 16035 473 16271
rect 709 16035 795 16271
rect 1031 16035 1117 16271
rect 1353 16035 1439 16271
rect 1675 16035 1761 16271
rect 1997 16035 2083 16271
rect 2319 16035 2405 16271
rect 2641 16035 2727 16271
rect 2963 16035 3049 16271
rect 3285 16035 3371 16271
rect 3607 16035 3693 16271
rect 3929 16035 4015 16271
rect 4251 16035 4337 16271
rect 4573 16035 4659 16271
rect 4895 16035 4981 16271
rect 5217 16035 5303 16271
rect 5539 16035 5830 16271
rect 8 15935 5830 16035
rect 8 15699 151 15935
rect 387 15699 473 15935
rect 709 15699 795 15935
rect 1031 15699 1117 15935
rect 1353 15699 1439 15935
rect 1675 15699 1761 15935
rect 1997 15699 2083 15935
rect 2319 15699 2405 15935
rect 2641 15699 2727 15935
rect 2963 15699 3049 15935
rect 3285 15699 3371 15935
rect 3607 15699 3693 15935
rect 3929 15699 4015 15935
rect 4251 15699 4337 15935
rect 4573 15699 4659 15935
rect 4895 15699 4981 15935
rect 5217 15699 5303 15935
rect 5539 15699 5830 15935
rect 8 15599 5830 15699
rect 8 15363 151 15599
rect 387 15363 473 15599
rect 709 15363 795 15599
rect 1031 15363 1117 15599
rect 1353 15363 1439 15599
rect 1675 15363 1761 15599
rect 1997 15363 2083 15599
rect 2319 15363 2405 15599
rect 2641 15363 2727 15599
rect 2963 15363 3049 15599
rect 3285 15363 3371 15599
rect 3607 15363 3693 15599
rect 3929 15363 4015 15599
rect 4251 15363 4337 15599
rect 4573 15363 4659 15599
rect 4895 15363 4981 15599
rect 5217 15363 5303 15599
rect 5539 15363 5830 15599
rect 8 15263 5830 15363
rect 8 15027 151 15263
rect 387 15027 473 15263
rect 709 15027 795 15263
rect 1031 15027 1117 15263
rect 1353 15027 1439 15263
rect 1675 15027 1761 15263
rect 1997 15027 2083 15263
rect 2319 15027 2405 15263
rect 2641 15027 2727 15263
rect 2963 15027 3049 15263
rect 3285 15027 3371 15263
rect 3607 15027 3693 15263
rect 3929 15027 4015 15263
rect 4251 15027 4337 15263
rect 4573 15027 4659 15263
rect 4895 15027 4981 15263
rect 5217 15027 5303 15263
rect 5539 15027 5830 15263
rect 8 14927 5830 15027
rect 8 14691 151 14927
rect 387 14691 473 14927
rect 709 14691 795 14927
rect 1031 14691 1117 14927
rect 1353 14691 1439 14927
rect 1675 14691 1761 14927
rect 1997 14691 2083 14927
rect 2319 14691 2405 14927
rect 2641 14691 2727 14927
rect 2963 14691 3049 14927
rect 3285 14691 3371 14927
rect 3607 14691 3693 14927
rect 3929 14691 4015 14927
rect 4251 14691 4337 14927
rect 4573 14691 4659 14927
rect 4895 14691 4981 14927
rect 5217 14691 5303 14927
rect 5539 14691 5830 14927
rect 8 14591 5830 14691
rect 8 14355 151 14591
rect 387 14355 473 14591
rect 709 14355 795 14591
rect 1031 14355 1117 14591
rect 1353 14355 1439 14591
rect 1675 14355 1761 14591
rect 1997 14355 2083 14591
rect 2319 14355 2405 14591
rect 2641 14355 2727 14591
rect 2963 14355 3049 14591
rect 3285 14355 3371 14591
rect 3607 14355 3693 14591
rect 3929 14355 4015 14591
rect 4251 14355 4337 14591
rect 4573 14355 4659 14591
rect 4895 14355 4981 14591
rect 5217 14355 5303 14591
rect 5539 14355 5830 14591
rect 8 14255 5830 14355
rect 8 14019 151 14255
rect 387 14019 473 14255
rect 709 14019 795 14255
rect 1031 14019 1117 14255
rect 1353 14019 1439 14255
rect 1675 14019 1761 14255
rect 1997 14019 2083 14255
rect 2319 14019 2405 14255
rect 2641 14019 2727 14255
rect 2963 14019 3049 14255
rect 3285 14019 3371 14255
rect 3607 14019 3693 14255
rect 3929 14019 4015 14255
rect 4251 14019 4337 14255
rect 4573 14019 4659 14255
rect 4895 14019 4981 14255
rect 5217 14019 5303 14255
rect 5539 14194 5830 14255
rect 5539 14019 5630 14194
rect 8 13994 5630 14019
tri 5630 13994 5830 14194 nw
tri 9148 18787 9348 18987 se
rect 9348 18959 15008 18987
rect 9348 18787 9477 18959
rect 9148 18723 9477 18787
rect 9713 18723 9798 18959
rect 10034 18723 10119 18959
rect 10355 18723 10440 18959
rect 10676 18723 10761 18959
rect 10997 18723 11082 18959
rect 11318 18723 11403 18959
rect 11639 18723 11724 18959
rect 11960 18723 12045 18959
rect 12281 18723 12366 18959
rect 12602 18723 12687 18959
rect 12923 18723 13008 18959
rect 13244 18723 13329 18959
rect 13565 18723 13650 18959
rect 13886 18723 13971 18959
rect 14207 18723 14292 18959
rect 14528 18723 14613 18959
rect 14849 18723 15008 18959
rect 9148 18623 15008 18723
rect 9148 18387 9477 18623
rect 9713 18387 9798 18623
rect 10034 18387 10119 18623
rect 10355 18387 10440 18623
rect 10676 18387 10761 18623
rect 10997 18387 11082 18623
rect 11318 18387 11403 18623
rect 11639 18387 11724 18623
rect 11960 18387 12045 18623
rect 12281 18387 12366 18623
rect 12602 18387 12687 18623
rect 12923 18387 13008 18623
rect 13244 18387 13329 18623
rect 13565 18387 13650 18623
rect 13886 18387 13971 18623
rect 14207 18387 14292 18623
rect 14528 18387 14613 18623
rect 14849 18387 15008 18623
rect 9148 18287 15008 18387
rect 9148 18051 9477 18287
rect 9713 18051 9798 18287
rect 10034 18051 10119 18287
rect 10355 18051 10440 18287
rect 10676 18051 10761 18287
rect 10997 18051 11082 18287
rect 11318 18051 11403 18287
rect 11639 18051 11724 18287
rect 11960 18051 12045 18287
rect 12281 18051 12366 18287
rect 12602 18051 12687 18287
rect 12923 18051 13008 18287
rect 13244 18051 13329 18287
rect 13565 18051 13650 18287
rect 13886 18051 13971 18287
rect 14207 18051 14292 18287
rect 14528 18051 14613 18287
rect 14849 18051 15008 18287
rect 9148 17951 15008 18051
rect 9148 17715 9477 17951
rect 9713 17715 9798 17951
rect 10034 17715 10119 17951
rect 10355 17715 10440 17951
rect 10676 17715 10761 17951
rect 10997 17715 11082 17951
rect 11318 17715 11403 17951
rect 11639 17715 11724 17951
rect 11960 17715 12045 17951
rect 12281 17715 12366 17951
rect 12602 17715 12687 17951
rect 12923 17715 13008 17951
rect 13244 17715 13329 17951
rect 13565 17715 13650 17951
rect 13886 17715 13971 17951
rect 14207 17715 14292 17951
rect 14528 17715 14613 17951
rect 14849 17715 15008 17951
rect 9148 17615 15008 17715
rect 9148 17379 9477 17615
rect 9713 17379 9798 17615
rect 10034 17379 10119 17615
rect 10355 17379 10440 17615
rect 10676 17379 10761 17615
rect 10997 17379 11082 17615
rect 11318 17379 11403 17615
rect 11639 17379 11724 17615
rect 11960 17379 12045 17615
rect 12281 17379 12366 17615
rect 12602 17379 12687 17615
rect 12923 17379 13008 17615
rect 13244 17379 13329 17615
rect 13565 17379 13650 17615
rect 13886 17379 13971 17615
rect 14207 17379 14292 17615
rect 14528 17379 14613 17615
rect 14849 17379 15008 17615
rect 9148 17279 15008 17379
rect 9148 17043 9477 17279
rect 9713 17043 9798 17279
rect 10034 17043 10119 17279
rect 10355 17043 10440 17279
rect 10676 17043 10761 17279
rect 10997 17043 11082 17279
rect 11318 17043 11403 17279
rect 11639 17043 11724 17279
rect 11960 17043 12045 17279
rect 12281 17043 12366 17279
rect 12602 17043 12687 17279
rect 12923 17043 13008 17279
rect 13244 17043 13329 17279
rect 13565 17043 13650 17279
rect 13886 17043 13971 17279
rect 14207 17043 14292 17279
rect 14528 17043 14613 17279
rect 14849 17043 15008 17279
rect 9148 16943 15008 17043
rect 9148 16707 9477 16943
rect 9713 16707 9798 16943
rect 10034 16707 10119 16943
rect 10355 16707 10440 16943
rect 10676 16707 10761 16943
rect 10997 16707 11082 16943
rect 11318 16707 11403 16943
rect 11639 16707 11724 16943
rect 11960 16707 12045 16943
rect 12281 16707 12366 16943
rect 12602 16707 12687 16943
rect 12923 16707 13008 16943
rect 13244 16707 13329 16943
rect 13565 16707 13650 16943
rect 13886 16707 13971 16943
rect 14207 16707 14292 16943
rect 14528 16707 14613 16943
rect 14849 16707 15008 16943
rect 9148 16607 15008 16707
rect 9148 16371 9477 16607
rect 9713 16371 9798 16607
rect 10034 16371 10119 16607
rect 10355 16371 10440 16607
rect 10676 16371 10761 16607
rect 10997 16371 11082 16607
rect 11318 16371 11403 16607
rect 11639 16371 11724 16607
rect 11960 16371 12045 16607
rect 12281 16371 12366 16607
rect 12602 16371 12687 16607
rect 12923 16371 13008 16607
rect 13244 16371 13329 16607
rect 13565 16371 13650 16607
rect 13886 16371 13971 16607
rect 14207 16371 14292 16607
rect 14528 16371 14613 16607
rect 14849 16371 15008 16607
rect 9148 16271 15008 16371
rect 9148 16035 9477 16271
rect 9713 16035 9798 16271
rect 10034 16035 10119 16271
rect 10355 16035 10440 16271
rect 10676 16035 10761 16271
rect 10997 16035 11082 16271
rect 11318 16035 11403 16271
rect 11639 16035 11724 16271
rect 11960 16035 12045 16271
rect 12281 16035 12366 16271
rect 12602 16035 12687 16271
rect 12923 16035 13008 16271
rect 13244 16035 13329 16271
rect 13565 16035 13650 16271
rect 13886 16035 13971 16271
rect 14207 16035 14292 16271
rect 14528 16035 14613 16271
rect 14849 16035 15008 16271
rect 9148 15935 15008 16035
rect 9148 15699 9477 15935
rect 9713 15699 9798 15935
rect 10034 15699 10119 15935
rect 10355 15699 10440 15935
rect 10676 15699 10761 15935
rect 10997 15699 11082 15935
rect 11318 15699 11403 15935
rect 11639 15699 11724 15935
rect 11960 15699 12045 15935
rect 12281 15699 12366 15935
rect 12602 15699 12687 15935
rect 12923 15699 13008 15935
rect 13244 15699 13329 15935
rect 13565 15699 13650 15935
rect 13886 15699 13971 15935
rect 14207 15699 14292 15935
rect 14528 15699 14613 15935
rect 14849 15699 15008 15935
rect 9148 15599 15008 15699
rect 9148 15363 9477 15599
rect 9713 15363 9798 15599
rect 10034 15363 10119 15599
rect 10355 15363 10440 15599
rect 10676 15363 10761 15599
rect 10997 15363 11082 15599
rect 11318 15363 11403 15599
rect 11639 15363 11724 15599
rect 11960 15363 12045 15599
rect 12281 15363 12366 15599
rect 12602 15363 12687 15599
rect 12923 15363 13008 15599
rect 13244 15363 13329 15599
rect 13565 15363 13650 15599
rect 13886 15363 13971 15599
rect 14207 15363 14292 15599
rect 14528 15363 14613 15599
rect 14849 15363 15008 15599
rect 9148 15263 15008 15363
rect 9148 15027 9477 15263
rect 9713 15027 9798 15263
rect 10034 15027 10119 15263
rect 10355 15027 10440 15263
rect 10676 15027 10761 15263
rect 10997 15027 11082 15263
rect 11318 15027 11403 15263
rect 11639 15027 11724 15263
rect 11960 15027 12045 15263
rect 12281 15027 12366 15263
rect 12602 15027 12687 15263
rect 12923 15027 13008 15263
rect 13244 15027 13329 15263
rect 13565 15027 13650 15263
rect 13886 15027 13971 15263
rect 14207 15027 14292 15263
rect 14528 15027 14613 15263
rect 14849 15027 15008 15263
rect 9148 14927 15008 15027
rect 9148 14691 9477 14927
rect 9713 14691 9798 14927
rect 10034 14691 10119 14927
rect 10355 14691 10440 14927
rect 10676 14691 10761 14927
rect 10997 14691 11082 14927
rect 11318 14691 11403 14927
rect 11639 14691 11724 14927
rect 11960 14691 12045 14927
rect 12281 14691 12366 14927
rect 12602 14691 12687 14927
rect 12923 14691 13008 14927
rect 13244 14691 13329 14927
rect 13565 14691 13650 14927
rect 13886 14691 13971 14927
rect 14207 14691 14292 14927
rect 14528 14691 14613 14927
rect 14849 14691 15008 14927
rect 9148 14591 15008 14691
rect 9148 14355 9477 14591
rect 9713 14355 9798 14591
rect 10034 14355 10119 14591
rect 10355 14355 10440 14591
rect 10676 14355 10761 14591
rect 10997 14355 11082 14591
rect 11318 14355 11403 14591
rect 11639 14355 11724 14591
rect 11960 14355 12045 14591
rect 12281 14355 12366 14591
rect 12602 14355 12687 14591
rect 12923 14355 13008 14591
rect 13244 14355 13329 14591
rect 13565 14355 13650 14591
rect 13886 14355 13971 14591
rect 14207 14355 14292 14591
rect 14528 14355 14613 14591
rect 14849 14355 15008 14591
rect 9148 14255 15008 14355
rect 9148 14194 9477 14255
tri 9148 13994 9348 14194 ne
rect 9348 14019 9477 14194
rect 9713 14019 9798 14255
rect 10034 14019 10119 14255
rect 10355 14019 10440 14255
rect 10676 14019 10761 14255
rect 10997 14019 11082 14255
rect 11318 14019 11403 14255
rect 11639 14019 11724 14255
rect 11960 14019 12045 14255
rect 12281 14019 12366 14255
rect 12602 14019 12687 14255
rect 12923 14019 13008 14255
rect 13244 14019 13329 14255
rect 13565 14019 13650 14255
rect 13886 14019 13971 14255
rect 14207 14019 14292 14255
rect 14528 14019 14613 14255
rect 14849 14019 15008 14255
rect 9348 13994 15008 14019
<< via4 >>
rect 249 39716 485 39952
rect 576 39716 812 39952
rect 903 39716 1139 39952
rect 1230 39716 1466 39952
rect 1557 39716 1793 39952
rect 1884 39716 2120 39952
rect 2211 39716 2447 39952
rect 2538 39716 2774 39952
rect 2865 39716 3101 39952
rect 3192 39716 3428 39952
rect 3519 39716 3755 39952
rect 3846 39716 4082 39952
rect 4173 39716 4409 39952
rect 4500 39716 4736 39952
rect 4827 39716 5063 39952
rect 5154 39716 5390 39952
rect 5481 39716 5717 39952
rect 5808 39716 6044 39952
rect 6135 39716 6371 39952
rect 6462 39716 6698 39952
rect 6789 39716 7025 39952
rect 7116 39716 7352 39952
rect 7443 39716 7679 39952
rect 7770 39716 8006 39952
rect 8097 39716 8333 39952
rect 8423 39716 8659 39952
rect 8749 39716 8985 39952
rect 9075 39716 9311 39952
rect 9401 39716 9637 39952
rect 9727 39716 9963 39952
rect 10053 39716 10289 39952
rect 10379 39716 10615 39952
rect 10705 39716 10941 39952
rect 11031 39716 11267 39952
rect 11357 39716 11593 39952
rect 11683 39716 11919 39952
rect 12009 39716 12245 39952
rect 12335 39716 12571 39952
rect 12661 39716 12897 39952
rect 12987 39716 13223 39952
rect 13313 39716 13549 39952
rect 13639 39716 13875 39952
rect 13965 39716 14201 39952
rect 14291 39716 14527 39952
rect 14617 39716 14853 39952
rect 249 39392 485 39628
rect 576 39392 812 39628
rect 903 39392 1139 39628
rect 1230 39392 1466 39628
rect 1557 39392 1793 39628
rect 1884 39392 2120 39628
rect 2211 39392 2447 39628
rect 2538 39392 2774 39628
rect 2865 39392 3101 39628
rect 3192 39392 3428 39628
rect 3519 39392 3755 39628
rect 3846 39392 4082 39628
rect 4173 39392 4409 39628
rect 4500 39392 4736 39628
rect 4827 39392 5063 39628
rect 5154 39392 5390 39628
rect 5481 39392 5717 39628
rect 5808 39392 6044 39628
rect 6135 39392 6371 39628
rect 6462 39392 6698 39628
rect 6789 39392 7025 39628
rect 7116 39392 7352 39628
rect 7443 39392 7679 39628
rect 7770 39392 8006 39628
rect 8097 39392 8333 39628
rect 8423 39392 8659 39628
rect 8749 39392 8985 39628
rect 9075 39392 9311 39628
rect 9401 39392 9637 39628
rect 9727 39392 9963 39628
rect 10053 39392 10289 39628
rect 10379 39392 10615 39628
rect 10705 39392 10941 39628
rect 11031 39392 11267 39628
rect 11357 39392 11593 39628
rect 11683 39392 11919 39628
rect 12009 39392 12245 39628
rect 12335 39392 12571 39628
rect 12661 39392 12897 39628
rect 12987 39392 13223 39628
rect 13313 39392 13549 39628
rect 13639 39392 13875 39628
rect 13965 39392 14201 39628
rect 14291 39392 14527 39628
rect 14617 39392 14853 39628
rect 249 39068 485 39304
rect 576 39068 812 39304
rect 903 39068 1139 39304
rect 1230 39068 1466 39304
rect 1557 39068 1793 39304
rect 1884 39068 2120 39304
rect 2211 39068 2447 39304
rect 2538 39068 2774 39304
rect 2865 39068 3101 39304
rect 3192 39068 3428 39304
rect 3519 39068 3755 39304
rect 3846 39068 4082 39304
rect 4173 39068 4409 39304
rect 4500 39068 4736 39304
rect 4827 39068 5063 39304
rect 5154 39068 5390 39304
rect 5481 39068 5717 39304
rect 5808 39068 6044 39304
rect 6135 39068 6371 39304
rect 6462 39068 6698 39304
rect 6789 39068 7025 39304
rect 7116 39068 7352 39304
rect 7443 39068 7679 39304
rect 7770 39068 8006 39304
rect 8097 39068 8333 39304
rect 8423 39068 8659 39304
rect 8749 39068 8985 39304
rect 9075 39068 9311 39304
rect 9401 39068 9637 39304
rect 9727 39068 9963 39304
rect 10053 39068 10289 39304
rect 10379 39068 10615 39304
rect 10705 39068 10941 39304
rect 11031 39068 11267 39304
rect 11357 39068 11593 39304
rect 11683 39068 11919 39304
rect 12009 39068 12245 39304
rect 12335 39068 12571 39304
rect 12661 39068 12897 39304
rect 12987 39068 13223 39304
rect 13313 39068 13549 39304
rect 13639 39068 13875 39304
rect 13965 39068 14201 39304
rect 14291 39068 14527 39304
rect 14617 39068 14853 39304
rect 249 38744 485 38980
rect 576 38744 812 38980
rect 903 38744 1139 38980
rect 1230 38744 1466 38980
rect 1557 38744 1793 38980
rect 1884 38744 2120 38980
rect 2211 38744 2447 38980
rect 2538 38744 2774 38980
rect 2865 38744 3101 38980
rect 3192 38744 3428 38980
rect 3519 38744 3755 38980
rect 3846 38744 4082 38980
rect 4173 38744 4409 38980
rect 4500 38744 4736 38980
rect 4827 38744 5063 38980
rect 5154 38744 5390 38980
rect 5481 38744 5717 38980
rect 5808 38744 6044 38980
rect 6135 38744 6371 38980
rect 6462 38744 6698 38980
rect 6789 38744 7025 38980
rect 7116 38744 7352 38980
rect 7443 38744 7679 38980
rect 7770 38744 8006 38980
rect 8097 38744 8333 38980
rect 8423 38744 8659 38980
rect 8749 38744 8985 38980
rect 9075 38744 9311 38980
rect 9401 38744 9637 38980
rect 9727 38744 9963 38980
rect 10053 38744 10289 38980
rect 10379 38744 10615 38980
rect 10705 38744 10941 38980
rect 11031 38744 11267 38980
rect 11357 38744 11593 38980
rect 11683 38744 11919 38980
rect 12009 38744 12245 38980
rect 12335 38744 12571 38980
rect 12661 38744 12897 38980
rect 12987 38744 13223 38980
rect 13313 38744 13549 38980
rect 13639 38744 13875 38980
rect 13965 38744 14201 38980
rect 14291 38744 14527 38980
rect 14617 38744 14853 38980
rect 249 38420 485 38656
rect 576 38420 812 38656
rect 903 38420 1139 38656
rect 1230 38420 1466 38656
rect 1557 38420 1793 38656
rect 1884 38420 2120 38656
rect 2211 38420 2447 38656
rect 2538 38420 2774 38656
rect 2865 38420 3101 38656
rect 3192 38420 3428 38656
rect 3519 38420 3755 38656
rect 3846 38420 4082 38656
rect 4173 38420 4409 38656
rect 4500 38420 4736 38656
rect 4827 38420 5063 38656
rect 5154 38420 5390 38656
rect 5481 38420 5717 38656
rect 5808 38420 6044 38656
rect 6135 38420 6371 38656
rect 6462 38420 6698 38656
rect 6789 38420 7025 38656
rect 7116 38420 7352 38656
rect 7443 38420 7679 38656
rect 7770 38420 8006 38656
rect 8097 38420 8333 38656
rect 8423 38420 8659 38656
rect 8749 38420 8985 38656
rect 9075 38420 9311 38656
rect 9401 38420 9637 38656
rect 9727 38420 9963 38656
rect 10053 38420 10289 38656
rect 10379 38420 10615 38656
rect 10705 38420 10941 38656
rect 11031 38420 11267 38656
rect 11357 38420 11593 38656
rect 11683 38420 11919 38656
rect 12009 38420 12245 38656
rect 12335 38420 12571 38656
rect 12661 38420 12897 38656
rect 12987 38420 13223 38656
rect 13313 38420 13549 38656
rect 13639 38420 13875 38656
rect 13965 38420 14201 38656
rect 14291 38420 14527 38656
rect 14617 38420 14853 38656
rect 249 38096 485 38332
rect 576 38096 812 38332
rect 903 38096 1139 38332
rect 1230 38096 1466 38332
rect 1557 38096 1793 38332
rect 1884 38096 2120 38332
rect 2211 38096 2447 38332
rect 2538 38096 2774 38332
rect 2865 38096 3101 38332
rect 3192 38096 3428 38332
rect 3519 38096 3755 38332
rect 3846 38096 4082 38332
rect 4173 38096 4409 38332
rect 4500 38096 4736 38332
rect 4827 38096 5063 38332
rect 5154 38096 5390 38332
rect 5481 38096 5717 38332
rect 5808 38096 6044 38332
rect 6135 38096 6371 38332
rect 6462 38096 6698 38332
rect 6789 38096 7025 38332
rect 7116 38096 7352 38332
rect 7443 38096 7679 38332
rect 7770 38096 8006 38332
rect 8097 38096 8333 38332
rect 8423 38096 8659 38332
rect 8749 38096 8985 38332
rect 9075 38096 9311 38332
rect 9401 38096 9637 38332
rect 9727 38096 9963 38332
rect 10053 38096 10289 38332
rect 10379 38096 10615 38332
rect 10705 38096 10941 38332
rect 11031 38096 11267 38332
rect 11357 38096 11593 38332
rect 11683 38096 11919 38332
rect 12009 38096 12245 38332
rect 12335 38096 12571 38332
rect 12661 38096 12897 38332
rect 12987 38096 13223 38332
rect 13313 38096 13549 38332
rect 13639 38096 13875 38332
rect 13965 38096 14201 38332
rect 14291 38096 14527 38332
rect 14617 38096 14853 38332
rect 249 37772 485 38008
rect 576 37772 812 38008
rect 903 37772 1139 38008
rect 1230 37772 1466 38008
rect 1557 37772 1793 38008
rect 1884 37772 2120 38008
rect 2211 37772 2447 38008
rect 2538 37772 2774 38008
rect 2865 37772 3101 38008
rect 3192 37772 3428 38008
rect 3519 37772 3755 38008
rect 3846 37772 4082 38008
rect 4173 37772 4409 38008
rect 4500 37772 4736 38008
rect 4827 37772 5063 38008
rect 5154 37772 5390 38008
rect 5481 37772 5717 38008
rect 5808 37772 6044 38008
rect 6135 37772 6371 38008
rect 6462 37772 6698 38008
rect 6789 37772 7025 38008
rect 7116 37772 7352 38008
rect 7443 37772 7679 38008
rect 7770 37772 8006 38008
rect 8097 37772 8333 38008
rect 8423 37772 8659 38008
rect 8749 37772 8985 38008
rect 9075 37772 9311 38008
rect 9401 37772 9637 38008
rect 9727 37772 9963 38008
rect 10053 37772 10289 38008
rect 10379 37772 10615 38008
rect 10705 37772 10941 38008
rect 11031 37772 11267 38008
rect 11357 37772 11593 38008
rect 11683 37772 11919 38008
rect 12009 37772 12245 38008
rect 12335 37772 12571 38008
rect 12661 37772 12897 38008
rect 12987 37772 13223 38008
rect 13313 37772 13549 38008
rect 13639 37772 13875 38008
rect 13965 37772 14201 38008
rect 14291 37772 14527 38008
rect 14617 37772 14853 38008
rect 249 37448 485 37684
rect 576 37448 812 37684
rect 903 37448 1139 37684
rect 1230 37448 1466 37684
rect 1557 37448 1793 37684
rect 1884 37448 2120 37684
rect 2211 37448 2447 37684
rect 2538 37448 2774 37684
rect 2865 37448 3101 37684
rect 3192 37448 3428 37684
rect 3519 37448 3755 37684
rect 3846 37448 4082 37684
rect 4173 37448 4409 37684
rect 4500 37448 4736 37684
rect 4827 37448 5063 37684
rect 5154 37448 5390 37684
rect 5481 37448 5717 37684
rect 5808 37448 6044 37684
rect 6135 37448 6371 37684
rect 6462 37448 6698 37684
rect 6789 37448 7025 37684
rect 7116 37448 7352 37684
rect 7443 37448 7679 37684
rect 7770 37448 8006 37684
rect 8097 37448 8333 37684
rect 8423 37448 8659 37684
rect 8749 37448 8985 37684
rect 9075 37448 9311 37684
rect 9401 37448 9637 37684
rect 9727 37448 9963 37684
rect 10053 37448 10289 37684
rect 10379 37448 10615 37684
rect 10705 37448 10941 37684
rect 11031 37448 11267 37684
rect 11357 37448 11593 37684
rect 11683 37448 11919 37684
rect 12009 37448 12245 37684
rect 12335 37448 12571 37684
rect 12661 37448 12897 37684
rect 12987 37448 13223 37684
rect 13313 37448 13549 37684
rect 13639 37448 13875 37684
rect 13965 37448 14201 37684
rect 14291 37448 14527 37684
rect 14617 37448 14853 37684
rect 249 37124 485 37360
rect 576 37124 812 37360
rect 903 37124 1139 37360
rect 1230 37124 1466 37360
rect 1557 37124 1793 37360
rect 1884 37124 2120 37360
rect 2211 37124 2447 37360
rect 2538 37124 2774 37360
rect 2865 37124 3101 37360
rect 3192 37124 3428 37360
rect 3519 37124 3755 37360
rect 3846 37124 4082 37360
rect 4173 37124 4409 37360
rect 4500 37124 4736 37360
rect 4827 37124 5063 37360
rect 5154 37124 5390 37360
rect 5481 37124 5717 37360
rect 5808 37124 6044 37360
rect 6135 37124 6371 37360
rect 6462 37124 6698 37360
rect 6789 37124 7025 37360
rect 7116 37124 7352 37360
rect 7443 37124 7679 37360
rect 7770 37124 8006 37360
rect 8097 37124 8333 37360
rect 8423 37124 8659 37360
rect 8749 37124 8985 37360
rect 9075 37124 9311 37360
rect 9401 37124 9637 37360
rect 9727 37124 9963 37360
rect 10053 37124 10289 37360
rect 10379 37124 10615 37360
rect 10705 37124 10941 37360
rect 11031 37124 11267 37360
rect 11357 37124 11593 37360
rect 11683 37124 11919 37360
rect 12009 37124 12245 37360
rect 12335 37124 12571 37360
rect 12661 37124 12897 37360
rect 12987 37124 13223 37360
rect 13313 37124 13549 37360
rect 13639 37124 13875 37360
rect 13965 37124 14201 37360
rect 14291 37124 14527 37360
rect 14617 37124 14853 37360
rect 249 36800 485 37036
rect 576 36800 812 37036
rect 903 36800 1139 37036
rect 1230 36800 1466 37036
rect 1557 36800 1793 37036
rect 1884 36800 2120 37036
rect 2211 36800 2447 37036
rect 2538 36800 2774 37036
rect 2865 36800 3101 37036
rect 3192 36800 3428 37036
rect 3519 36800 3755 37036
rect 3846 36800 4082 37036
rect 4173 36800 4409 37036
rect 4500 36800 4736 37036
rect 4827 36800 5063 37036
rect 5154 36800 5390 37036
rect 5481 36800 5717 37036
rect 5808 36800 6044 37036
rect 6135 36800 6371 37036
rect 6462 36800 6698 37036
rect 6789 36800 7025 37036
rect 7116 36800 7352 37036
rect 7443 36800 7679 37036
rect 7770 36800 8006 37036
rect 8097 36800 8333 37036
rect 8423 36800 8659 37036
rect 8749 36800 8985 37036
rect 9075 36800 9311 37036
rect 9401 36800 9637 37036
rect 9727 36800 9963 37036
rect 10053 36800 10289 37036
rect 10379 36800 10615 37036
rect 10705 36800 10941 37036
rect 11031 36800 11267 37036
rect 11357 36800 11593 37036
rect 11683 36800 11919 37036
rect 12009 36800 12245 37036
rect 12335 36800 12571 37036
rect 12661 36800 12897 37036
rect 12987 36800 13223 37036
rect 13313 36800 13549 37036
rect 13639 36800 13875 37036
rect 13965 36800 14201 37036
rect 14291 36800 14527 37036
rect 14617 36800 14853 37036
rect 249 36476 485 36712
rect 576 36476 812 36712
rect 903 36476 1139 36712
rect 1230 36476 1466 36712
rect 1557 36476 1793 36712
rect 1884 36476 2120 36712
rect 2211 36476 2447 36712
rect 2538 36476 2774 36712
rect 2865 36476 3101 36712
rect 3192 36476 3428 36712
rect 3519 36476 3755 36712
rect 3846 36476 4082 36712
rect 4173 36476 4409 36712
rect 4500 36476 4736 36712
rect 4827 36476 5063 36712
rect 5154 36476 5390 36712
rect 5481 36476 5717 36712
rect 5808 36476 6044 36712
rect 6135 36476 6371 36712
rect 6462 36476 6698 36712
rect 6789 36476 7025 36712
rect 7116 36476 7352 36712
rect 7443 36476 7679 36712
rect 7770 36476 8006 36712
rect 8097 36476 8333 36712
rect 8423 36476 8659 36712
rect 8749 36476 8985 36712
rect 9075 36476 9311 36712
rect 9401 36476 9637 36712
rect 9727 36476 9963 36712
rect 10053 36476 10289 36712
rect 10379 36476 10615 36712
rect 10705 36476 10941 36712
rect 11031 36476 11267 36712
rect 11357 36476 11593 36712
rect 11683 36476 11919 36712
rect 12009 36476 12245 36712
rect 12335 36476 12571 36712
rect 12661 36476 12897 36712
rect 12987 36476 13223 36712
rect 13313 36476 13549 36712
rect 13639 36476 13875 36712
rect 13965 36476 14201 36712
rect 14291 36476 14527 36712
rect 14617 36476 14853 36712
rect 249 36152 485 36388
rect 576 36152 812 36388
rect 903 36152 1139 36388
rect 1230 36152 1466 36388
rect 1557 36152 1793 36388
rect 1884 36152 2120 36388
rect 2211 36152 2447 36388
rect 2538 36152 2774 36388
rect 2865 36152 3101 36388
rect 3192 36152 3428 36388
rect 3519 36152 3755 36388
rect 3846 36152 4082 36388
rect 4173 36152 4409 36388
rect 4500 36152 4736 36388
rect 4827 36152 5063 36388
rect 5154 36152 5390 36388
rect 5481 36152 5717 36388
rect 5808 36152 6044 36388
rect 6135 36152 6371 36388
rect 6462 36152 6698 36388
rect 6789 36152 7025 36388
rect 7116 36152 7352 36388
rect 7443 36152 7679 36388
rect 7770 36152 8006 36388
rect 8097 36152 8333 36388
rect 8423 36152 8659 36388
rect 8749 36152 8985 36388
rect 9075 36152 9311 36388
rect 9401 36152 9637 36388
rect 9727 36152 9963 36388
rect 10053 36152 10289 36388
rect 10379 36152 10615 36388
rect 10705 36152 10941 36388
rect 11031 36152 11267 36388
rect 11357 36152 11593 36388
rect 11683 36152 11919 36388
rect 12009 36152 12245 36388
rect 12335 36152 12571 36388
rect 12661 36152 12897 36388
rect 12987 36152 13223 36388
rect 13313 36152 13549 36388
rect 13639 36152 13875 36388
rect 13965 36152 14201 36388
rect 14291 36152 14527 36388
rect 14617 36152 14853 36388
rect 249 35828 485 36064
rect 576 35828 812 36064
rect 903 35828 1139 36064
rect 1230 35828 1466 36064
rect 1557 35828 1793 36064
rect 1884 35828 2120 36064
rect 2211 35828 2447 36064
rect 2538 35828 2774 36064
rect 2865 35828 3101 36064
rect 3192 35828 3428 36064
rect 3519 35828 3755 36064
rect 3846 35828 4082 36064
rect 4173 35828 4409 36064
rect 4500 35828 4736 36064
rect 4827 35828 5063 36064
rect 5154 35828 5390 36064
rect 5481 35828 5717 36064
rect 5808 35828 6044 36064
rect 6135 35828 6371 36064
rect 6462 35828 6698 36064
rect 6789 35828 7025 36064
rect 7116 35828 7352 36064
rect 7443 35828 7679 36064
rect 7770 35828 8006 36064
rect 8097 35828 8333 36064
rect 8423 35828 8659 36064
rect 8749 35828 8985 36064
rect 9075 35828 9311 36064
rect 9401 35828 9637 36064
rect 9727 35828 9963 36064
rect 10053 35828 10289 36064
rect 10379 35828 10615 36064
rect 10705 35828 10941 36064
rect 11031 35828 11267 36064
rect 11357 35828 11593 36064
rect 11683 35828 11919 36064
rect 12009 35828 12245 36064
rect 12335 35828 12571 36064
rect 12661 35828 12897 36064
rect 12987 35828 13223 36064
rect 13313 35828 13549 36064
rect 13639 35828 13875 36064
rect 13965 35828 14201 36064
rect 14291 35828 14527 36064
rect 14617 35828 14853 36064
rect 249 35504 485 35740
rect 576 35504 812 35740
rect 903 35504 1139 35740
rect 1230 35504 1466 35740
rect 1557 35504 1793 35740
rect 1884 35504 2120 35740
rect 2211 35504 2447 35740
rect 2538 35504 2774 35740
rect 2865 35504 3101 35740
rect 3192 35504 3428 35740
rect 3519 35504 3755 35740
rect 3846 35504 4082 35740
rect 4173 35504 4409 35740
rect 4500 35504 4736 35740
rect 4827 35504 5063 35740
rect 5154 35504 5390 35740
rect 5481 35504 5717 35740
rect 5808 35504 6044 35740
rect 6135 35504 6371 35740
rect 6462 35504 6698 35740
rect 6789 35504 7025 35740
rect 7116 35504 7352 35740
rect 7443 35504 7679 35740
rect 7770 35504 8006 35740
rect 8097 35504 8333 35740
rect 8423 35504 8659 35740
rect 8749 35504 8985 35740
rect 9075 35504 9311 35740
rect 9401 35504 9637 35740
rect 9727 35504 9963 35740
rect 10053 35504 10289 35740
rect 10379 35504 10615 35740
rect 10705 35504 10941 35740
rect 11031 35504 11267 35740
rect 11357 35504 11593 35740
rect 11683 35504 11919 35740
rect 12009 35504 12245 35740
rect 12335 35504 12571 35740
rect 12661 35504 12897 35740
rect 12987 35504 13223 35740
rect 13313 35504 13549 35740
rect 13639 35504 13875 35740
rect 13965 35504 14201 35740
rect 14291 35504 14527 35740
rect 14617 35504 14853 35740
rect 249 35180 485 35416
rect 576 35180 812 35416
rect 903 35180 1139 35416
rect 1230 35180 1466 35416
rect 1557 35180 1793 35416
rect 1884 35180 2120 35416
rect 2211 35180 2447 35416
rect 2538 35180 2774 35416
rect 2865 35180 3101 35416
rect 3192 35180 3428 35416
rect 3519 35180 3755 35416
rect 3846 35180 4082 35416
rect 4173 35180 4409 35416
rect 4500 35180 4736 35416
rect 4827 35180 5063 35416
rect 5154 35180 5390 35416
rect 5481 35180 5717 35416
rect 5808 35180 6044 35416
rect 6135 35180 6371 35416
rect 6462 35180 6698 35416
rect 6789 35180 7025 35416
rect 7116 35180 7352 35416
rect 7443 35180 7679 35416
rect 7770 35180 8006 35416
rect 8097 35180 8333 35416
rect 8423 35180 8659 35416
rect 8749 35180 8985 35416
rect 9075 35180 9311 35416
rect 9401 35180 9637 35416
rect 9727 35180 9963 35416
rect 10053 35180 10289 35416
rect 10379 35180 10615 35416
rect 10705 35180 10941 35416
rect 11031 35180 11267 35416
rect 11357 35180 11593 35416
rect 11683 35180 11919 35416
rect 12009 35180 12245 35416
rect 12335 35180 12571 35416
rect 12661 35180 12897 35416
rect 12987 35180 13223 35416
rect 13313 35180 13549 35416
rect 13639 35180 13875 35416
rect 13965 35180 14201 35416
rect 14291 35180 14527 35416
rect 14617 35180 14853 35416
rect 151 18723 387 18959
rect 473 18723 709 18959
rect 795 18723 1031 18959
rect 1117 18723 1353 18959
rect 1439 18723 1675 18959
rect 1761 18723 1997 18959
rect 2083 18723 2319 18959
rect 2405 18723 2641 18959
rect 2727 18723 2963 18959
rect 3049 18723 3285 18959
rect 3371 18723 3607 18959
rect 3693 18723 3929 18959
rect 4015 18723 4251 18959
rect 4337 18723 4573 18959
rect 4659 18723 4895 18959
rect 4981 18723 5217 18959
rect 5303 18723 5539 18959
rect 151 18387 387 18623
rect 473 18387 709 18623
rect 795 18387 1031 18623
rect 1117 18387 1353 18623
rect 1439 18387 1675 18623
rect 1761 18387 1997 18623
rect 2083 18387 2319 18623
rect 2405 18387 2641 18623
rect 2727 18387 2963 18623
rect 3049 18387 3285 18623
rect 3371 18387 3607 18623
rect 3693 18387 3929 18623
rect 4015 18387 4251 18623
rect 4337 18387 4573 18623
rect 4659 18387 4895 18623
rect 4981 18387 5217 18623
rect 5303 18387 5539 18623
rect 151 18051 387 18287
rect 473 18051 709 18287
rect 795 18051 1031 18287
rect 1117 18051 1353 18287
rect 1439 18051 1675 18287
rect 1761 18051 1997 18287
rect 2083 18051 2319 18287
rect 2405 18051 2641 18287
rect 2727 18051 2963 18287
rect 3049 18051 3285 18287
rect 3371 18051 3607 18287
rect 3693 18051 3929 18287
rect 4015 18051 4251 18287
rect 4337 18051 4573 18287
rect 4659 18051 4895 18287
rect 4981 18051 5217 18287
rect 5303 18051 5539 18287
rect 151 17715 387 17951
rect 473 17715 709 17951
rect 795 17715 1031 17951
rect 1117 17715 1353 17951
rect 1439 17715 1675 17951
rect 1761 17715 1997 17951
rect 2083 17715 2319 17951
rect 2405 17715 2641 17951
rect 2727 17715 2963 17951
rect 3049 17715 3285 17951
rect 3371 17715 3607 17951
rect 3693 17715 3929 17951
rect 4015 17715 4251 17951
rect 4337 17715 4573 17951
rect 4659 17715 4895 17951
rect 4981 17715 5217 17951
rect 5303 17715 5539 17951
rect 151 17379 387 17615
rect 473 17379 709 17615
rect 795 17379 1031 17615
rect 1117 17379 1353 17615
rect 1439 17379 1675 17615
rect 1761 17379 1997 17615
rect 2083 17379 2319 17615
rect 2405 17379 2641 17615
rect 2727 17379 2963 17615
rect 3049 17379 3285 17615
rect 3371 17379 3607 17615
rect 3693 17379 3929 17615
rect 4015 17379 4251 17615
rect 4337 17379 4573 17615
rect 4659 17379 4895 17615
rect 4981 17379 5217 17615
rect 5303 17379 5539 17615
rect 151 17043 387 17279
rect 473 17043 709 17279
rect 795 17043 1031 17279
rect 1117 17043 1353 17279
rect 1439 17043 1675 17279
rect 1761 17043 1997 17279
rect 2083 17043 2319 17279
rect 2405 17043 2641 17279
rect 2727 17043 2963 17279
rect 3049 17043 3285 17279
rect 3371 17043 3607 17279
rect 3693 17043 3929 17279
rect 4015 17043 4251 17279
rect 4337 17043 4573 17279
rect 4659 17043 4895 17279
rect 4981 17043 5217 17279
rect 5303 17043 5539 17279
rect 151 16707 387 16943
rect 473 16707 709 16943
rect 795 16707 1031 16943
rect 1117 16707 1353 16943
rect 1439 16707 1675 16943
rect 1761 16707 1997 16943
rect 2083 16707 2319 16943
rect 2405 16707 2641 16943
rect 2727 16707 2963 16943
rect 3049 16707 3285 16943
rect 3371 16707 3607 16943
rect 3693 16707 3929 16943
rect 4015 16707 4251 16943
rect 4337 16707 4573 16943
rect 4659 16707 4895 16943
rect 4981 16707 5217 16943
rect 5303 16707 5539 16943
rect 151 16371 387 16607
rect 473 16371 709 16607
rect 795 16371 1031 16607
rect 1117 16371 1353 16607
rect 1439 16371 1675 16607
rect 1761 16371 1997 16607
rect 2083 16371 2319 16607
rect 2405 16371 2641 16607
rect 2727 16371 2963 16607
rect 3049 16371 3285 16607
rect 3371 16371 3607 16607
rect 3693 16371 3929 16607
rect 4015 16371 4251 16607
rect 4337 16371 4573 16607
rect 4659 16371 4895 16607
rect 4981 16371 5217 16607
rect 5303 16371 5539 16607
rect 151 16035 387 16271
rect 473 16035 709 16271
rect 795 16035 1031 16271
rect 1117 16035 1353 16271
rect 1439 16035 1675 16271
rect 1761 16035 1997 16271
rect 2083 16035 2319 16271
rect 2405 16035 2641 16271
rect 2727 16035 2963 16271
rect 3049 16035 3285 16271
rect 3371 16035 3607 16271
rect 3693 16035 3929 16271
rect 4015 16035 4251 16271
rect 4337 16035 4573 16271
rect 4659 16035 4895 16271
rect 4981 16035 5217 16271
rect 5303 16035 5539 16271
rect 151 15699 387 15935
rect 473 15699 709 15935
rect 795 15699 1031 15935
rect 1117 15699 1353 15935
rect 1439 15699 1675 15935
rect 1761 15699 1997 15935
rect 2083 15699 2319 15935
rect 2405 15699 2641 15935
rect 2727 15699 2963 15935
rect 3049 15699 3285 15935
rect 3371 15699 3607 15935
rect 3693 15699 3929 15935
rect 4015 15699 4251 15935
rect 4337 15699 4573 15935
rect 4659 15699 4895 15935
rect 4981 15699 5217 15935
rect 5303 15699 5539 15935
rect 151 15363 387 15599
rect 473 15363 709 15599
rect 795 15363 1031 15599
rect 1117 15363 1353 15599
rect 1439 15363 1675 15599
rect 1761 15363 1997 15599
rect 2083 15363 2319 15599
rect 2405 15363 2641 15599
rect 2727 15363 2963 15599
rect 3049 15363 3285 15599
rect 3371 15363 3607 15599
rect 3693 15363 3929 15599
rect 4015 15363 4251 15599
rect 4337 15363 4573 15599
rect 4659 15363 4895 15599
rect 4981 15363 5217 15599
rect 5303 15363 5539 15599
rect 151 15027 387 15263
rect 473 15027 709 15263
rect 795 15027 1031 15263
rect 1117 15027 1353 15263
rect 1439 15027 1675 15263
rect 1761 15027 1997 15263
rect 2083 15027 2319 15263
rect 2405 15027 2641 15263
rect 2727 15027 2963 15263
rect 3049 15027 3285 15263
rect 3371 15027 3607 15263
rect 3693 15027 3929 15263
rect 4015 15027 4251 15263
rect 4337 15027 4573 15263
rect 4659 15027 4895 15263
rect 4981 15027 5217 15263
rect 5303 15027 5539 15263
rect 151 14691 387 14927
rect 473 14691 709 14927
rect 795 14691 1031 14927
rect 1117 14691 1353 14927
rect 1439 14691 1675 14927
rect 1761 14691 1997 14927
rect 2083 14691 2319 14927
rect 2405 14691 2641 14927
rect 2727 14691 2963 14927
rect 3049 14691 3285 14927
rect 3371 14691 3607 14927
rect 3693 14691 3929 14927
rect 4015 14691 4251 14927
rect 4337 14691 4573 14927
rect 4659 14691 4895 14927
rect 4981 14691 5217 14927
rect 5303 14691 5539 14927
rect 151 14355 387 14591
rect 473 14355 709 14591
rect 795 14355 1031 14591
rect 1117 14355 1353 14591
rect 1439 14355 1675 14591
rect 1761 14355 1997 14591
rect 2083 14355 2319 14591
rect 2405 14355 2641 14591
rect 2727 14355 2963 14591
rect 3049 14355 3285 14591
rect 3371 14355 3607 14591
rect 3693 14355 3929 14591
rect 4015 14355 4251 14591
rect 4337 14355 4573 14591
rect 4659 14355 4895 14591
rect 4981 14355 5217 14591
rect 5303 14355 5539 14591
rect 151 14019 387 14255
rect 473 14019 709 14255
rect 795 14019 1031 14255
rect 1117 14019 1353 14255
rect 1439 14019 1675 14255
rect 1761 14019 1997 14255
rect 2083 14019 2319 14255
rect 2405 14019 2641 14255
rect 2727 14019 2963 14255
rect 3049 14019 3285 14255
rect 3371 14019 3607 14255
rect 3693 14019 3929 14255
rect 4015 14019 4251 14255
rect 4337 14019 4573 14255
rect 4659 14019 4895 14255
rect 4981 14019 5217 14255
rect 5303 14019 5539 14255
rect 9477 18723 9713 18959
rect 9798 18723 10034 18959
rect 10119 18723 10355 18959
rect 10440 18723 10676 18959
rect 10761 18723 10997 18959
rect 11082 18723 11318 18959
rect 11403 18723 11639 18959
rect 11724 18723 11960 18959
rect 12045 18723 12281 18959
rect 12366 18723 12602 18959
rect 12687 18723 12923 18959
rect 13008 18723 13244 18959
rect 13329 18723 13565 18959
rect 13650 18723 13886 18959
rect 13971 18723 14207 18959
rect 14292 18723 14528 18959
rect 14613 18723 14849 18959
rect 9477 18387 9713 18623
rect 9798 18387 10034 18623
rect 10119 18387 10355 18623
rect 10440 18387 10676 18623
rect 10761 18387 10997 18623
rect 11082 18387 11318 18623
rect 11403 18387 11639 18623
rect 11724 18387 11960 18623
rect 12045 18387 12281 18623
rect 12366 18387 12602 18623
rect 12687 18387 12923 18623
rect 13008 18387 13244 18623
rect 13329 18387 13565 18623
rect 13650 18387 13886 18623
rect 13971 18387 14207 18623
rect 14292 18387 14528 18623
rect 14613 18387 14849 18623
rect 9477 18051 9713 18287
rect 9798 18051 10034 18287
rect 10119 18051 10355 18287
rect 10440 18051 10676 18287
rect 10761 18051 10997 18287
rect 11082 18051 11318 18287
rect 11403 18051 11639 18287
rect 11724 18051 11960 18287
rect 12045 18051 12281 18287
rect 12366 18051 12602 18287
rect 12687 18051 12923 18287
rect 13008 18051 13244 18287
rect 13329 18051 13565 18287
rect 13650 18051 13886 18287
rect 13971 18051 14207 18287
rect 14292 18051 14528 18287
rect 14613 18051 14849 18287
rect 9477 17715 9713 17951
rect 9798 17715 10034 17951
rect 10119 17715 10355 17951
rect 10440 17715 10676 17951
rect 10761 17715 10997 17951
rect 11082 17715 11318 17951
rect 11403 17715 11639 17951
rect 11724 17715 11960 17951
rect 12045 17715 12281 17951
rect 12366 17715 12602 17951
rect 12687 17715 12923 17951
rect 13008 17715 13244 17951
rect 13329 17715 13565 17951
rect 13650 17715 13886 17951
rect 13971 17715 14207 17951
rect 14292 17715 14528 17951
rect 14613 17715 14849 17951
rect 9477 17379 9713 17615
rect 9798 17379 10034 17615
rect 10119 17379 10355 17615
rect 10440 17379 10676 17615
rect 10761 17379 10997 17615
rect 11082 17379 11318 17615
rect 11403 17379 11639 17615
rect 11724 17379 11960 17615
rect 12045 17379 12281 17615
rect 12366 17379 12602 17615
rect 12687 17379 12923 17615
rect 13008 17379 13244 17615
rect 13329 17379 13565 17615
rect 13650 17379 13886 17615
rect 13971 17379 14207 17615
rect 14292 17379 14528 17615
rect 14613 17379 14849 17615
rect 9477 17043 9713 17279
rect 9798 17043 10034 17279
rect 10119 17043 10355 17279
rect 10440 17043 10676 17279
rect 10761 17043 10997 17279
rect 11082 17043 11318 17279
rect 11403 17043 11639 17279
rect 11724 17043 11960 17279
rect 12045 17043 12281 17279
rect 12366 17043 12602 17279
rect 12687 17043 12923 17279
rect 13008 17043 13244 17279
rect 13329 17043 13565 17279
rect 13650 17043 13886 17279
rect 13971 17043 14207 17279
rect 14292 17043 14528 17279
rect 14613 17043 14849 17279
rect 9477 16707 9713 16943
rect 9798 16707 10034 16943
rect 10119 16707 10355 16943
rect 10440 16707 10676 16943
rect 10761 16707 10997 16943
rect 11082 16707 11318 16943
rect 11403 16707 11639 16943
rect 11724 16707 11960 16943
rect 12045 16707 12281 16943
rect 12366 16707 12602 16943
rect 12687 16707 12923 16943
rect 13008 16707 13244 16943
rect 13329 16707 13565 16943
rect 13650 16707 13886 16943
rect 13971 16707 14207 16943
rect 14292 16707 14528 16943
rect 14613 16707 14849 16943
rect 9477 16371 9713 16607
rect 9798 16371 10034 16607
rect 10119 16371 10355 16607
rect 10440 16371 10676 16607
rect 10761 16371 10997 16607
rect 11082 16371 11318 16607
rect 11403 16371 11639 16607
rect 11724 16371 11960 16607
rect 12045 16371 12281 16607
rect 12366 16371 12602 16607
rect 12687 16371 12923 16607
rect 13008 16371 13244 16607
rect 13329 16371 13565 16607
rect 13650 16371 13886 16607
rect 13971 16371 14207 16607
rect 14292 16371 14528 16607
rect 14613 16371 14849 16607
rect 9477 16035 9713 16271
rect 9798 16035 10034 16271
rect 10119 16035 10355 16271
rect 10440 16035 10676 16271
rect 10761 16035 10997 16271
rect 11082 16035 11318 16271
rect 11403 16035 11639 16271
rect 11724 16035 11960 16271
rect 12045 16035 12281 16271
rect 12366 16035 12602 16271
rect 12687 16035 12923 16271
rect 13008 16035 13244 16271
rect 13329 16035 13565 16271
rect 13650 16035 13886 16271
rect 13971 16035 14207 16271
rect 14292 16035 14528 16271
rect 14613 16035 14849 16271
rect 9477 15699 9713 15935
rect 9798 15699 10034 15935
rect 10119 15699 10355 15935
rect 10440 15699 10676 15935
rect 10761 15699 10997 15935
rect 11082 15699 11318 15935
rect 11403 15699 11639 15935
rect 11724 15699 11960 15935
rect 12045 15699 12281 15935
rect 12366 15699 12602 15935
rect 12687 15699 12923 15935
rect 13008 15699 13244 15935
rect 13329 15699 13565 15935
rect 13650 15699 13886 15935
rect 13971 15699 14207 15935
rect 14292 15699 14528 15935
rect 14613 15699 14849 15935
rect 9477 15363 9713 15599
rect 9798 15363 10034 15599
rect 10119 15363 10355 15599
rect 10440 15363 10676 15599
rect 10761 15363 10997 15599
rect 11082 15363 11318 15599
rect 11403 15363 11639 15599
rect 11724 15363 11960 15599
rect 12045 15363 12281 15599
rect 12366 15363 12602 15599
rect 12687 15363 12923 15599
rect 13008 15363 13244 15599
rect 13329 15363 13565 15599
rect 13650 15363 13886 15599
rect 13971 15363 14207 15599
rect 14292 15363 14528 15599
rect 14613 15363 14849 15599
rect 9477 15027 9713 15263
rect 9798 15027 10034 15263
rect 10119 15027 10355 15263
rect 10440 15027 10676 15263
rect 10761 15027 10997 15263
rect 11082 15027 11318 15263
rect 11403 15027 11639 15263
rect 11724 15027 11960 15263
rect 12045 15027 12281 15263
rect 12366 15027 12602 15263
rect 12687 15027 12923 15263
rect 13008 15027 13244 15263
rect 13329 15027 13565 15263
rect 13650 15027 13886 15263
rect 13971 15027 14207 15263
rect 14292 15027 14528 15263
rect 14613 15027 14849 15263
rect 9477 14691 9713 14927
rect 9798 14691 10034 14927
rect 10119 14691 10355 14927
rect 10440 14691 10676 14927
rect 10761 14691 10997 14927
rect 11082 14691 11318 14927
rect 11403 14691 11639 14927
rect 11724 14691 11960 14927
rect 12045 14691 12281 14927
rect 12366 14691 12602 14927
rect 12687 14691 12923 14927
rect 13008 14691 13244 14927
rect 13329 14691 13565 14927
rect 13650 14691 13886 14927
rect 13971 14691 14207 14927
rect 14292 14691 14528 14927
rect 14613 14691 14849 14927
rect 9477 14355 9713 14591
rect 9798 14355 10034 14591
rect 10119 14355 10355 14591
rect 10440 14355 10676 14591
rect 10761 14355 10997 14591
rect 11082 14355 11318 14591
rect 11403 14355 11639 14591
rect 11724 14355 11960 14591
rect 12045 14355 12281 14591
rect 12366 14355 12602 14591
rect 12687 14355 12923 14591
rect 13008 14355 13244 14591
rect 13329 14355 13565 14591
rect 13650 14355 13886 14591
rect 13971 14355 14207 14591
rect 14292 14355 14528 14591
rect 14613 14355 14849 14591
rect 9477 14019 9713 14255
rect 9798 14019 10034 14255
rect 10119 14019 10355 14255
rect 10440 14019 10676 14255
rect 10761 14019 10997 14255
rect 11082 14019 11318 14255
rect 11403 14019 11639 14255
rect 11724 14019 11960 14255
rect 12045 14019 12281 14255
rect 12366 14019 12602 14255
rect 12687 14019 12923 14255
rect 13008 14019 13244 14255
rect 13329 14019 13565 14255
rect 13650 14019 13886 14255
rect 13971 14019 14207 14255
rect 14292 14019 14528 14255
rect 14613 14019 14849 14255
<< metal5 >>
rect 8 39952 15008 39987
rect 8 39716 249 39952
rect 485 39716 576 39952
rect 812 39716 903 39952
rect 1139 39716 1230 39952
rect 1466 39716 1557 39952
rect 1793 39716 1884 39952
rect 2120 39716 2211 39952
rect 2447 39716 2538 39952
rect 2774 39716 2865 39952
rect 3101 39716 3192 39952
rect 3428 39716 3519 39952
rect 3755 39716 3846 39952
rect 4082 39716 4173 39952
rect 4409 39716 4500 39952
rect 4736 39716 4827 39952
rect 5063 39716 5154 39952
rect 5390 39716 5481 39952
rect 5717 39716 5808 39952
rect 6044 39716 6135 39952
rect 6371 39716 6462 39952
rect 6698 39716 6789 39952
rect 7025 39716 7116 39952
rect 7352 39716 7443 39952
rect 7679 39716 7770 39952
rect 8006 39716 8097 39952
rect 8333 39716 8423 39952
rect 8659 39716 8749 39952
rect 8985 39716 9075 39952
rect 9311 39716 9401 39952
rect 9637 39716 9727 39952
rect 9963 39716 10053 39952
rect 10289 39716 10379 39952
rect 10615 39716 10705 39952
rect 10941 39716 11031 39952
rect 11267 39716 11357 39952
rect 11593 39716 11683 39952
rect 11919 39716 12009 39952
rect 12245 39716 12335 39952
rect 12571 39716 12661 39952
rect 12897 39716 12987 39952
rect 13223 39716 13313 39952
rect 13549 39716 13639 39952
rect 13875 39716 13965 39952
rect 14201 39716 14291 39952
rect 14527 39716 14617 39952
rect 14853 39716 15008 39952
rect 8 39628 15008 39716
rect 8 39392 249 39628
rect 485 39392 576 39628
rect 812 39392 903 39628
rect 1139 39392 1230 39628
rect 1466 39392 1557 39628
rect 1793 39392 1884 39628
rect 2120 39392 2211 39628
rect 2447 39392 2538 39628
rect 2774 39392 2865 39628
rect 3101 39392 3192 39628
rect 3428 39392 3519 39628
rect 3755 39392 3846 39628
rect 4082 39392 4173 39628
rect 4409 39392 4500 39628
rect 4736 39392 4827 39628
rect 5063 39392 5154 39628
rect 5390 39392 5481 39628
rect 5717 39392 5808 39628
rect 6044 39392 6135 39628
rect 6371 39392 6462 39628
rect 6698 39392 6789 39628
rect 7025 39392 7116 39628
rect 7352 39392 7443 39628
rect 7679 39392 7770 39628
rect 8006 39392 8097 39628
rect 8333 39392 8423 39628
rect 8659 39392 8749 39628
rect 8985 39392 9075 39628
rect 9311 39392 9401 39628
rect 9637 39392 9727 39628
rect 9963 39392 10053 39628
rect 10289 39392 10379 39628
rect 10615 39392 10705 39628
rect 10941 39392 11031 39628
rect 11267 39392 11357 39628
rect 11593 39392 11683 39628
rect 11919 39392 12009 39628
rect 12245 39392 12335 39628
rect 12571 39392 12661 39628
rect 12897 39392 12987 39628
rect 13223 39392 13313 39628
rect 13549 39392 13639 39628
rect 13875 39392 13965 39628
rect 14201 39392 14291 39628
rect 14527 39392 14617 39628
rect 14853 39392 15008 39628
rect 8 39304 15008 39392
rect 8 39068 249 39304
rect 485 39068 576 39304
rect 812 39068 903 39304
rect 1139 39068 1230 39304
rect 1466 39068 1557 39304
rect 1793 39068 1884 39304
rect 2120 39068 2211 39304
rect 2447 39068 2538 39304
rect 2774 39068 2865 39304
rect 3101 39068 3192 39304
rect 3428 39068 3519 39304
rect 3755 39068 3846 39304
rect 4082 39068 4173 39304
rect 4409 39068 4500 39304
rect 4736 39068 4827 39304
rect 5063 39068 5154 39304
rect 5390 39068 5481 39304
rect 5717 39068 5808 39304
rect 6044 39068 6135 39304
rect 6371 39068 6462 39304
rect 6698 39068 6789 39304
rect 7025 39068 7116 39304
rect 7352 39068 7443 39304
rect 7679 39068 7770 39304
rect 8006 39068 8097 39304
rect 8333 39068 8423 39304
rect 8659 39068 8749 39304
rect 8985 39068 9075 39304
rect 9311 39068 9401 39304
rect 9637 39068 9727 39304
rect 9963 39068 10053 39304
rect 10289 39068 10379 39304
rect 10615 39068 10705 39304
rect 10941 39068 11031 39304
rect 11267 39068 11357 39304
rect 11593 39068 11683 39304
rect 11919 39068 12009 39304
rect 12245 39068 12335 39304
rect 12571 39068 12661 39304
rect 12897 39068 12987 39304
rect 13223 39068 13313 39304
rect 13549 39068 13639 39304
rect 13875 39068 13965 39304
rect 14201 39068 14291 39304
rect 14527 39068 14617 39304
rect 14853 39068 15008 39304
rect 8 38980 15008 39068
rect 8 38744 249 38980
rect 485 38744 576 38980
rect 812 38744 903 38980
rect 1139 38744 1230 38980
rect 1466 38744 1557 38980
rect 1793 38744 1884 38980
rect 2120 38744 2211 38980
rect 2447 38744 2538 38980
rect 2774 38744 2865 38980
rect 3101 38744 3192 38980
rect 3428 38744 3519 38980
rect 3755 38744 3846 38980
rect 4082 38744 4173 38980
rect 4409 38744 4500 38980
rect 4736 38744 4827 38980
rect 5063 38744 5154 38980
rect 5390 38744 5481 38980
rect 5717 38744 5808 38980
rect 6044 38744 6135 38980
rect 6371 38744 6462 38980
rect 6698 38744 6789 38980
rect 7025 38744 7116 38980
rect 7352 38744 7443 38980
rect 7679 38744 7770 38980
rect 8006 38744 8097 38980
rect 8333 38744 8423 38980
rect 8659 38744 8749 38980
rect 8985 38744 9075 38980
rect 9311 38744 9401 38980
rect 9637 38744 9727 38980
rect 9963 38744 10053 38980
rect 10289 38744 10379 38980
rect 10615 38744 10705 38980
rect 10941 38744 11031 38980
rect 11267 38744 11357 38980
rect 11593 38744 11683 38980
rect 11919 38744 12009 38980
rect 12245 38744 12335 38980
rect 12571 38744 12661 38980
rect 12897 38744 12987 38980
rect 13223 38744 13313 38980
rect 13549 38744 13639 38980
rect 13875 38744 13965 38980
rect 14201 38744 14291 38980
rect 14527 38744 14617 38980
rect 14853 38744 15008 38980
rect 8 38656 15008 38744
rect 8 38420 249 38656
rect 485 38420 576 38656
rect 812 38420 903 38656
rect 1139 38420 1230 38656
rect 1466 38420 1557 38656
rect 1793 38420 1884 38656
rect 2120 38420 2211 38656
rect 2447 38420 2538 38656
rect 2774 38420 2865 38656
rect 3101 38420 3192 38656
rect 3428 38420 3519 38656
rect 3755 38420 3846 38656
rect 4082 38420 4173 38656
rect 4409 38420 4500 38656
rect 4736 38420 4827 38656
rect 5063 38420 5154 38656
rect 5390 38420 5481 38656
rect 5717 38420 5808 38656
rect 6044 38420 6135 38656
rect 6371 38420 6462 38656
rect 6698 38420 6789 38656
rect 7025 38420 7116 38656
rect 7352 38420 7443 38656
rect 7679 38420 7770 38656
rect 8006 38420 8097 38656
rect 8333 38420 8423 38656
rect 8659 38420 8749 38656
rect 8985 38420 9075 38656
rect 9311 38420 9401 38656
rect 9637 38420 9727 38656
rect 9963 38420 10053 38656
rect 10289 38420 10379 38656
rect 10615 38420 10705 38656
rect 10941 38420 11031 38656
rect 11267 38420 11357 38656
rect 11593 38420 11683 38656
rect 11919 38420 12009 38656
rect 12245 38420 12335 38656
rect 12571 38420 12661 38656
rect 12897 38420 12987 38656
rect 13223 38420 13313 38656
rect 13549 38420 13639 38656
rect 13875 38420 13965 38656
rect 14201 38420 14291 38656
rect 14527 38420 14617 38656
rect 14853 38420 15008 38656
rect 8 38332 15008 38420
rect 8 38096 249 38332
rect 485 38096 576 38332
rect 812 38096 903 38332
rect 1139 38096 1230 38332
rect 1466 38096 1557 38332
rect 1793 38096 1884 38332
rect 2120 38096 2211 38332
rect 2447 38096 2538 38332
rect 2774 38096 2865 38332
rect 3101 38096 3192 38332
rect 3428 38096 3519 38332
rect 3755 38096 3846 38332
rect 4082 38096 4173 38332
rect 4409 38096 4500 38332
rect 4736 38096 4827 38332
rect 5063 38096 5154 38332
rect 5390 38096 5481 38332
rect 5717 38096 5808 38332
rect 6044 38096 6135 38332
rect 6371 38096 6462 38332
rect 6698 38096 6789 38332
rect 7025 38096 7116 38332
rect 7352 38096 7443 38332
rect 7679 38096 7770 38332
rect 8006 38096 8097 38332
rect 8333 38096 8423 38332
rect 8659 38096 8749 38332
rect 8985 38096 9075 38332
rect 9311 38096 9401 38332
rect 9637 38096 9727 38332
rect 9963 38096 10053 38332
rect 10289 38096 10379 38332
rect 10615 38096 10705 38332
rect 10941 38096 11031 38332
rect 11267 38096 11357 38332
rect 11593 38096 11683 38332
rect 11919 38096 12009 38332
rect 12245 38096 12335 38332
rect 12571 38096 12661 38332
rect 12897 38096 12987 38332
rect 13223 38096 13313 38332
rect 13549 38096 13639 38332
rect 13875 38096 13965 38332
rect 14201 38096 14291 38332
rect 14527 38096 14617 38332
rect 14853 38096 15008 38332
rect 8 38008 15008 38096
rect 8 37772 249 38008
rect 485 37772 576 38008
rect 812 37772 903 38008
rect 1139 37772 1230 38008
rect 1466 37772 1557 38008
rect 1793 37772 1884 38008
rect 2120 37772 2211 38008
rect 2447 37772 2538 38008
rect 2774 37772 2865 38008
rect 3101 37772 3192 38008
rect 3428 37772 3519 38008
rect 3755 37772 3846 38008
rect 4082 37772 4173 38008
rect 4409 37772 4500 38008
rect 4736 37772 4827 38008
rect 5063 37772 5154 38008
rect 5390 37772 5481 38008
rect 5717 37772 5808 38008
rect 6044 37772 6135 38008
rect 6371 37772 6462 38008
rect 6698 37772 6789 38008
rect 7025 37772 7116 38008
rect 7352 37772 7443 38008
rect 7679 37772 7770 38008
rect 8006 37772 8097 38008
rect 8333 37772 8423 38008
rect 8659 37772 8749 38008
rect 8985 37772 9075 38008
rect 9311 37772 9401 38008
rect 9637 37772 9727 38008
rect 9963 37772 10053 38008
rect 10289 37772 10379 38008
rect 10615 37772 10705 38008
rect 10941 37772 11031 38008
rect 11267 37772 11357 38008
rect 11593 37772 11683 38008
rect 11919 37772 12009 38008
rect 12245 37772 12335 38008
rect 12571 37772 12661 38008
rect 12897 37772 12987 38008
rect 13223 37772 13313 38008
rect 13549 37772 13639 38008
rect 13875 37772 13965 38008
rect 14201 37772 14291 38008
rect 14527 37772 14617 38008
rect 14853 37772 15008 38008
rect 8 37684 15008 37772
rect 8 37448 249 37684
rect 485 37448 576 37684
rect 812 37448 903 37684
rect 1139 37448 1230 37684
rect 1466 37448 1557 37684
rect 1793 37448 1884 37684
rect 2120 37448 2211 37684
rect 2447 37448 2538 37684
rect 2774 37448 2865 37684
rect 3101 37448 3192 37684
rect 3428 37448 3519 37684
rect 3755 37448 3846 37684
rect 4082 37448 4173 37684
rect 4409 37448 4500 37684
rect 4736 37448 4827 37684
rect 5063 37448 5154 37684
rect 5390 37448 5481 37684
rect 5717 37448 5808 37684
rect 6044 37448 6135 37684
rect 6371 37448 6462 37684
rect 6698 37448 6789 37684
rect 7025 37448 7116 37684
rect 7352 37448 7443 37684
rect 7679 37448 7770 37684
rect 8006 37448 8097 37684
rect 8333 37448 8423 37684
rect 8659 37448 8749 37684
rect 8985 37448 9075 37684
rect 9311 37448 9401 37684
rect 9637 37448 9727 37684
rect 9963 37448 10053 37684
rect 10289 37448 10379 37684
rect 10615 37448 10705 37684
rect 10941 37448 11031 37684
rect 11267 37448 11357 37684
rect 11593 37448 11683 37684
rect 11919 37448 12009 37684
rect 12245 37448 12335 37684
rect 12571 37448 12661 37684
rect 12897 37448 12987 37684
rect 13223 37448 13313 37684
rect 13549 37448 13639 37684
rect 13875 37448 13965 37684
rect 14201 37448 14291 37684
rect 14527 37448 14617 37684
rect 14853 37448 15008 37684
rect 8 37360 15008 37448
rect 8 37124 249 37360
rect 485 37124 576 37360
rect 812 37124 903 37360
rect 1139 37124 1230 37360
rect 1466 37124 1557 37360
rect 1793 37124 1884 37360
rect 2120 37124 2211 37360
rect 2447 37124 2538 37360
rect 2774 37124 2865 37360
rect 3101 37124 3192 37360
rect 3428 37124 3519 37360
rect 3755 37124 3846 37360
rect 4082 37124 4173 37360
rect 4409 37124 4500 37360
rect 4736 37124 4827 37360
rect 5063 37124 5154 37360
rect 5390 37124 5481 37360
rect 5717 37124 5808 37360
rect 6044 37124 6135 37360
rect 6371 37124 6462 37360
rect 6698 37124 6789 37360
rect 7025 37124 7116 37360
rect 7352 37124 7443 37360
rect 7679 37124 7770 37360
rect 8006 37124 8097 37360
rect 8333 37124 8423 37360
rect 8659 37124 8749 37360
rect 8985 37124 9075 37360
rect 9311 37124 9401 37360
rect 9637 37124 9727 37360
rect 9963 37124 10053 37360
rect 10289 37124 10379 37360
rect 10615 37124 10705 37360
rect 10941 37124 11031 37360
rect 11267 37124 11357 37360
rect 11593 37124 11683 37360
rect 11919 37124 12009 37360
rect 12245 37124 12335 37360
rect 12571 37124 12661 37360
rect 12897 37124 12987 37360
rect 13223 37124 13313 37360
rect 13549 37124 13639 37360
rect 13875 37124 13965 37360
rect 14201 37124 14291 37360
rect 14527 37124 14617 37360
rect 14853 37124 15008 37360
rect 8 37036 15008 37124
rect 8 36800 249 37036
rect 485 36800 576 37036
rect 812 36800 903 37036
rect 1139 36800 1230 37036
rect 1466 36800 1557 37036
rect 1793 36800 1884 37036
rect 2120 36800 2211 37036
rect 2447 36800 2538 37036
rect 2774 36800 2865 37036
rect 3101 36800 3192 37036
rect 3428 36800 3519 37036
rect 3755 36800 3846 37036
rect 4082 36800 4173 37036
rect 4409 36800 4500 37036
rect 4736 36800 4827 37036
rect 5063 36800 5154 37036
rect 5390 36800 5481 37036
rect 5717 36800 5808 37036
rect 6044 36800 6135 37036
rect 6371 36800 6462 37036
rect 6698 36800 6789 37036
rect 7025 36800 7116 37036
rect 7352 36800 7443 37036
rect 7679 36800 7770 37036
rect 8006 36800 8097 37036
rect 8333 36800 8423 37036
rect 8659 36800 8749 37036
rect 8985 36800 9075 37036
rect 9311 36800 9401 37036
rect 9637 36800 9727 37036
rect 9963 36800 10053 37036
rect 10289 36800 10379 37036
rect 10615 36800 10705 37036
rect 10941 36800 11031 37036
rect 11267 36800 11357 37036
rect 11593 36800 11683 37036
rect 11919 36800 12009 37036
rect 12245 36800 12335 37036
rect 12571 36800 12661 37036
rect 12897 36800 12987 37036
rect 13223 36800 13313 37036
rect 13549 36800 13639 37036
rect 13875 36800 13965 37036
rect 14201 36800 14291 37036
rect 14527 36800 14617 37036
rect 14853 36800 15008 37036
rect 8 36712 15008 36800
rect 8 36476 249 36712
rect 485 36476 576 36712
rect 812 36476 903 36712
rect 1139 36476 1230 36712
rect 1466 36476 1557 36712
rect 1793 36476 1884 36712
rect 2120 36476 2211 36712
rect 2447 36476 2538 36712
rect 2774 36476 2865 36712
rect 3101 36476 3192 36712
rect 3428 36476 3519 36712
rect 3755 36476 3846 36712
rect 4082 36476 4173 36712
rect 4409 36476 4500 36712
rect 4736 36476 4827 36712
rect 5063 36476 5154 36712
rect 5390 36476 5481 36712
rect 5717 36476 5808 36712
rect 6044 36476 6135 36712
rect 6371 36476 6462 36712
rect 6698 36476 6789 36712
rect 7025 36476 7116 36712
rect 7352 36476 7443 36712
rect 7679 36476 7770 36712
rect 8006 36476 8097 36712
rect 8333 36476 8423 36712
rect 8659 36476 8749 36712
rect 8985 36476 9075 36712
rect 9311 36476 9401 36712
rect 9637 36476 9727 36712
rect 9963 36476 10053 36712
rect 10289 36476 10379 36712
rect 10615 36476 10705 36712
rect 10941 36476 11031 36712
rect 11267 36476 11357 36712
rect 11593 36476 11683 36712
rect 11919 36476 12009 36712
rect 12245 36476 12335 36712
rect 12571 36476 12661 36712
rect 12897 36476 12987 36712
rect 13223 36476 13313 36712
rect 13549 36476 13639 36712
rect 13875 36476 13965 36712
rect 14201 36476 14291 36712
rect 14527 36476 14617 36712
rect 14853 36476 15008 36712
rect 8 36388 15008 36476
rect 8 36152 249 36388
rect 485 36152 576 36388
rect 812 36152 903 36388
rect 1139 36152 1230 36388
rect 1466 36152 1557 36388
rect 1793 36152 1884 36388
rect 2120 36152 2211 36388
rect 2447 36152 2538 36388
rect 2774 36152 2865 36388
rect 3101 36152 3192 36388
rect 3428 36152 3519 36388
rect 3755 36152 3846 36388
rect 4082 36152 4173 36388
rect 4409 36152 4500 36388
rect 4736 36152 4827 36388
rect 5063 36152 5154 36388
rect 5390 36152 5481 36388
rect 5717 36152 5808 36388
rect 6044 36152 6135 36388
rect 6371 36152 6462 36388
rect 6698 36152 6789 36388
rect 7025 36152 7116 36388
rect 7352 36152 7443 36388
rect 7679 36152 7770 36388
rect 8006 36152 8097 36388
rect 8333 36152 8423 36388
rect 8659 36152 8749 36388
rect 8985 36152 9075 36388
rect 9311 36152 9401 36388
rect 9637 36152 9727 36388
rect 9963 36152 10053 36388
rect 10289 36152 10379 36388
rect 10615 36152 10705 36388
rect 10941 36152 11031 36388
rect 11267 36152 11357 36388
rect 11593 36152 11683 36388
rect 11919 36152 12009 36388
rect 12245 36152 12335 36388
rect 12571 36152 12661 36388
rect 12897 36152 12987 36388
rect 13223 36152 13313 36388
rect 13549 36152 13639 36388
rect 13875 36152 13965 36388
rect 14201 36152 14291 36388
rect 14527 36152 14617 36388
rect 14853 36152 15008 36388
rect 8 36064 15008 36152
rect 8 35828 249 36064
rect 485 35828 576 36064
rect 812 35828 903 36064
rect 1139 35828 1230 36064
rect 1466 35828 1557 36064
rect 1793 35828 1884 36064
rect 2120 35828 2211 36064
rect 2447 35828 2538 36064
rect 2774 35828 2865 36064
rect 3101 35828 3192 36064
rect 3428 35828 3519 36064
rect 3755 35828 3846 36064
rect 4082 35828 4173 36064
rect 4409 35828 4500 36064
rect 4736 35828 4827 36064
rect 5063 35828 5154 36064
rect 5390 35828 5481 36064
rect 5717 35828 5808 36064
rect 6044 35828 6135 36064
rect 6371 35828 6462 36064
rect 6698 35828 6789 36064
rect 7025 35828 7116 36064
rect 7352 35828 7443 36064
rect 7679 35828 7770 36064
rect 8006 35828 8097 36064
rect 8333 35828 8423 36064
rect 8659 35828 8749 36064
rect 8985 35828 9075 36064
rect 9311 35828 9401 36064
rect 9637 35828 9727 36064
rect 9963 35828 10053 36064
rect 10289 35828 10379 36064
rect 10615 35828 10705 36064
rect 10941 35828 11031 36064
rect 11267 35828 11357 36064
rect 11593 35828 11683 36064
rect 11919 35828 12009 36064
rect 12245 35828 12335 36064
rect 12571 35828 12661 36064
rect 12897 35828 12987 36064
rect 13223 35828 13313 36064
rect 13549 35828 13639 36064
rect 13875 35828 13965 36064
rect 14201 35828 14291 36064
rect 14527 35828 14617 36064
rect 14853 35828 15008 36064
rect 8 35740 15008 35828
rect 8 35504 249 35740
rect 485 35504 576 35740
rect 812 35504 903 35740
rect 1139 35504 1230 35740
rect 1466 35504 1557 35740
rect 1793 35504 1884 35740
rect 2120 35504 2211 35740
rect 2447 35504 2538 35740
rect 2774 35504 2865 35740
rect 3101 35504 3192 35740
rect 3428 35504 3519 35740
rect 3755 35504 3846 35740
rect 4082 35504 4173 35740
rect 4409 35504 4500 35740
rect 4736 35504 4827 35740
rect 5063 35504 5154 35740
rect 5390 35504 5481 35740
rect 5717 35504 5808 35740
rect 6044 35504 6135 35740
rect 6371 35504 6462 35740
rect 6698 35504 6789 35740
rect 7025 35504 7116 35740
rect 7352 35504 7443 35740
rect 7679 35504 7770 35740
rect 8006 35504 8097 35740
rect 8333 35504 8423 35740
rect 8659 35504 8749 35740
rect 8985 35504 9075 35740
rect 9311 35504 9401 35740
rect 9637 35504 9727 35740
rect 9963 35504 10053 35740
rect 10289 35504 10379 35740
rect 10615 35504 10705 35740
rect 10941 35504 11031 35740
rect 11267 35504 11357 35740
rect 11593 35504 11683 35740
rect 11919 35504 12009 35740
rect 12245 35504 12335 35740
rect 12571 35504 12661 35740
rect 12897 35504 12987 35740
rect 13223 35504 13313 35740
rect 13549 35504 13639 35740
rect 13875 35504 13965 35740
rect 14201 35504 14291 35740
rect 14527 35504 14617 35740
rect 14853 35504 15008 35740
rect 8 35416 15008 35504
rect 8 35180 249 35416
rect 485 35180 576 35416
rect 812 35180 903 35416
rect 1139 35180 1230 35416
rect 1466 35180 1557 35416
rect 1793 35180 1884 35416
rect 2120 35180 2211 35416
rect 2447 35180 2538 35416
rect 2774 35180 2865 35416
rect 3101 35180 3192 35416
rect 3428 35180 3519 35416
rect 3755 35180 3846 35416
rect 4082 35180 4173 35416
rect 4409 35180 4500 35416
rect 4736 35180 4827 35416
rect 5063 35180 5154 35416
rect 5390 35180 5481 35416
rect 5717 35180 5808 35416
rect 6044 35180 6135 35416
rect 6371 35180 6462 35416
rect 6698 35180 6789 35416
rect 7025 35180 7116 35416
rect 7352 35180 7443 35416
rect 7679 35180 7770 35416
rect 8006 35180 8097 35416
rect 8333 35180 8423 35416
rect 8659 35180 8749 35416
rect 8985 35180 9075 35416
rect 9311 35180 9401 35416
rect 9637 35180 9727 35416
rect 9963 35180 10053 35416
rect 10289 35180 10379 35416
rect 10615 35180 10705 35416
rect 10941 35180 11031 35416
rect 11267 35180 11357 35416
rect 11593 35180 11683 35416
rect 11919 35180 12009 35416
rect 12245 35180 12335 35416
rect 12571 35180 12661 35416
rect 12897 35180 12987 35416
rect 13223 35180 13313 35416
rect 13549 35180 13639 35416
rect 13875 35180 13965 35416
rect 14201 35180 14291 35416
rect 14527 35180 14617 35416
rect 14853 35180 15008 35416
rect 8 35144 15008 35180
rect 8 18959 15008 18984
rect 8 18723 151 18959
rect 387 18723 473 18959
rect 709 18723 795 18959
rect 1031 18723 1117 18959
rect 1353 18723 1439 18959
rect 1675 18723 1761 18959
rect 1997 18723 2083 18959
rect 2319 18723 2405 18959
rect 2641 18723 2727 18959
rect 2963 18723 3049 18959
rect 3285 18723 3371 18959
rect 3607 18723 3693 18959
rect 3929 18723 4015 18959
rect 4251 18723 4337 18959
rect 4573 18723 4659 18959
rect 4895 18723 4981 18959
rect 5217 18723 5303 18959
rect 5539 18723 9477 18959
rect 9713 18723 9798 18959
rect 10034 18723 10119 18959
rect 10355 18723 10440 18959
rect 10676 18723 10761 18959
rect 10997 18723 11082 18959
rect 11318 18723 11403 18959
rect 11639 18723 11724 18959
rect 11960 18723 12045 18959
rect 12281 18723 12366 18959
rect 12602 18723 12687 18959
rect 12923 18723 13008 18959
rect 13244 18723 13329 18959
rect 13565 18723 13650 18959
rect 13886 18723 13971 18959
rect 14207 18723 14292 18959
rect 14528 18723 14613 18959
rect 14849 18723 15008 18959
rect 8 18623 15008 18723
rect 8 18387 151 18623
rect 387 18387 473 18623
rect 709 18387 795 18623
rect 1031 18387 1117 18623
rect 1353 18387 1439 18623
rect 1675 18387 1761 18623
rect 1997 18387 2083 18623
rect 2319 18387 2405 18623
rect 2641 18387 2727 18623
rect 2963 18387 3049 18623
rect 3285 18387 3371 18623
rect 3607 18387 3693 18623
rect 3929 18387 4015 18623
rect 4251 18387 4337 18623
rect 4573 18387 4659 18623
rect 4895 18387 4981 18623
rect 5217 18387 5303 18623
rect 5539 18387 9477 18623
rect 9713 18387 9798 18623
rect 10034 18387 10119 18623
rect 10355 18387 10440 18623
rect 10676 18387 10761 18623
rect 10997 18387 11082 18623
rect 11318 18387 11403 18623
rect 11639 18387 11724 18623
rect 11960 18387 12045 18623
rect 12281 18387 12366 18623
rect 12602 18387 12687 18623
rect 12923 18387 13008 18623
rect 13244 18387 13329 18623
rect 13565 18387 13650 18623
rect 13886 18387 13971 18623
rect 14207 18387 14292 18623
rect 14528 18387 14613 18623
rect 14849 18387 15008 18623
rect 8 18287 15008 18387
rect 8 18051 151 18287
rect 387 18051 473 18287
rect 709 18051 795 18287
rect 1031 18051 1117 18287
rect 1353 18051 1439 18287
rect 1675 18051 1761 18287
rect 1997 18051 2083 18287
rect 2319 18051 2405 18287
rect 2641 18051 2727 18287
rect 2963 18051 3049 18287
rect 3285 18051 3371 18287
rect 3607 18051 3693 18287
rect 3929 18051 4015 18287
rect 4251 18051 4337 18287
rect 4573 18051 4659 18287
rect 4895 18051 4981 18287
rect 5217 18051 5303 18287
rect 5539 18051 9477 18287
rect 9713 18051 9798 18287
rect 10034 18051 10119 18287
rect 10355 18051 10440 18287
rect 10676 18051 10761 18287
rect 10997 18051 11082 18287
rect 11318 18051 11403 18287
rect 11639 18051 11724 18287
rect 11960 18051 12045 18287
rect 12281 18051 12366 18287
rect 12602 18051 12687 18287
rect 12923 18051 13008 18287
rect 13244 18051 13329 18287
rect 13565 18051 13650 18287
rect 13886 18051 13971 18287
rect 14207 18051 14292 18287
rect 14528 18051 14613 18287
rect 14849 18051 15008 18287
rect 8 17951 15008 18051
rect 8 17715 151 17951
rect 387 17715 473 17951
rect 709 17715 795 17951
rect 1031 17715 1117 17951
rect 1353 17715 1439 17951
rect 1675 17715 1761 17951
rect 1997 17715 2083 17951
rect 2319 17715 2405 17951
rect 2641 17715 2727 17951
rect 2963 17715 3049 17951
rect 3285 17715 3371 17951
rect 3607 17715 3693 17951
rect 3929 17715 4015 17951
rect 4251 17715 4337 17951
rect 4573 17715 4659 17951
rect 4895 17715 4981 17951
rect 5217 17715 5303 17951
rect 5539 17715 9477 17951
rect 9713 17715 9798 17951
rect 10034 17715 10119 17951
rect 10355 17715 10440 17951
rect 10676 17715 10761 17951
rect 10997 17715 11082 17951
rect 11318 17715 11403 17951
rect 11639 17715 11724 17951
rect 11960 17715 12045 17951
rect 12281 17715 12366 17951
rect 12602 17715 12687 17951
rect 12923 17715 13008 17951
rect 13244 17715 13329 17951
rect 13565 17715 13650 17951
rect 13886 17715 13971 17951
rect 14207 17715 14292 17951
rect 14528 17715 14613 17951
rect 14849 17715 15008 17951
rect 8 17615 15008 17715
rect 8 17379 151 17615
rect 387 17379 473 17615
rect 709 17379 795 17615
rect 1031 17379 1117 17615
rect 1353 17379 1439 17615
rect 1675 17379 1761 17615
rect 1997 17379 2083 17615
rect 2319 17379 2405 17615
rect 2641 17379 2727 17615
rect 2963 17379 3049 17615
rect 3285 17379 3371 17615
rect 3607 17379 3693 17615
rect 3929 17379 4015 17615
rect 4251 17379 4337 17615
rect 4573 17379 4659 17615
rect 4895 17379 4981 17615
rect 5217 17379 5303 17615
rect 5539 17379 9477 17615
rect 9713 17379 9798 17615
rect 10034 17379 10119 17615
rect 10355 17379 10440 17615
rect 10676 17379 10761 17615
rect 10997 17379 11082 17615
rect 11318 17379 11403 17615
rect 11639 17379 11724 17615
rect 11960 17379 12045 17615
rect 12281 17379 12366 17615
rect 12602 17379 12687 17615
rect 12923 17379 13008 17615
rect 13244 17379 13329 17615
rect 13565 17379 13650 17615
rect 13886 17379 13971 17615
rect 14207 17379 14292 17615
rect 14528 17379 14613 17615
rect 14849 17379 15008 17615
rect 8 17279 15008 17379
rect 8 17043 151 17279
rect 387 17043 473 17279
rect 709 17043 795 17279
rect 1031 17043 1117 17279
rect 1353 17043 1439 17279
rect 1675 17043 1761 17279
rect 1997 17043 2083 17279
rect 2319 17043 2405 17279
rect 2641 17043 2727 17279
rect 2963 17043 3049 17279
rect 3285 17043 3371 17279
rect 3607 17043 3693 17279
rect 3929 17043 4015 17279
rect 4251 17043 4337 17279
rect 4573 17043 4659 17279
rect 4895 17043 4981 17279
rect 5217 17043 5303 17279
rect 5539 17043 9477 17279
rect 9713 17043 9798 17279
rect 10034 17043 10119 17279
rect 10355 17043 10440 17279
rect 10676 17043 10761 17279
rect 10997 17043 11082 17279
rect 11318 17043 11403 17279
rect 11639 17043 11724 17279
rect 11960 17043 12045 17279
rect 12281 17043 12366 17279
rect 12602 17043 12687 17279
rect 12923 17043 13008 17279
rect 13244 17043 13329 17279
rect 13565 17043 13650 17279
rect 13886 17043 13971 17279
rect 14207 17043 14292 17279
rect 14528 17043 14613 17279
rect 14849 17043 15008 17279
rect 8 16943 15008 17043
rect 8 16707 151 16943
rect 387 16707 473 16943
rect 709 16707 795 16943
rect 1031 16707 1117 16943
rect 1353 16707 1439 16943
rect 1675 16707 1761 16943
rect 1997 16707 2083 16943
rect 2319 16707 2405 16943
rect 2641 16707 2727 16943
rect 2963 16707 3049 16943
rect 3285 16707 3371 16943
rect 3607 16707 3693 16943
rect 3929 16707 4015 16943
rect 4251 16707 4337 16943
rect 4573 16707 4659 16943
rect 4895 16707 4981 16943
rect 5217 16707 5303 16943
rect 5539 16707 9477 16943
rect 9713 16707 9798 16943
rect 10034 16707 10119 16943
rect 10355 16707 10440 16943
rect 10676 16707 10761 16943
rect 10997 16707 11082 16943
rect 11318 16707 11403 16943
rect 11639 16707 11724 16943
rect 11960 16707 12045 16943
rect 12281 16707 12366 16943
rect 12602 16707 12687 16943
rect 12923 16707 13008 16943
rect 13244 16707 13329 16943
rect 13565 16707 13650 16943
rect 13886 16707 13971 16943
rect 14207 16707 14292 16943
rect 14528 16707 14613 16943
rect 14849 16707 15008 16943
rect 8 16607 15008 16707
rect 8 16371 151 16607
rect 387 16371 473 16607
rect 709 16371 795 16607
rect 1031 16371 1117 16607
rect 1353 16371 1439 16607
rect 1675 16371 1761 16607
rect 1997 16371 2083 16607
rect 2319 16371 2405 16607
rect 2641 16371 2727 16607
rect 2963 16371 3049 16607
rect 3285 16371 3371 16607
rect 3607 16371 3693 16607
rect 3929 16371 4015 16607
rect 4251 16371 4337 16607
rect 4573 16371 4659 16607
rect 4895 16371 4981 16607
rect 5217 16371 5303 16607
rect 5539 16371 9477 16607
rect 9713 16371 9798 16607
rect 10034 16371 10119 16607
rect 10355 16371 10440 16607
rect 10676 16371 10761 16607
rect 10997 16371 11082 16607
rect 11318 16371 11403 16607
rect 11639 16371 11724 16607
rect 11960 16371 12045 16607
rect 12281 16371 12366 16607
rect 12602 16371 12687 16607
rect 12923 16371 13008 16607
rect 13244 16371 13329 16607
rect 13565 16371 13650 16607
rect 13886 16371 13971 16607
rect 14207 16371 14292 16607
rect 14528 16371 14613 16607
rect 14849 16371 15008 16607
rect 8 16271 15008 16371
rect 8 16035 151 16271
rect 387 16035 473 16271
rect 709 16035 795 16271
rect 1031 16035 1117 16271
rect 1353 16035 1439 16271
rect 1675 16035 1761 16271
rect 1997 16035 2083 16271
rect 2319 16035 2405 16271
rect 2641 16035 2727 16271
rect 2963 16035 3049 16271
rect 3285 16035 3371 16271
rect 3607 16035 3693 16271
rect 3929 16035 4015 16271
rect 4251 16035 4337 16271
rect 4573 16035 4659 16271
rect 4895 16035 4981 16271
rect 5217 16035 5303 16271
rect 5539 16035 9477 16271
rect 9713 16035 9798 16271
rect 10034 16035 10119 16271
rect 10355 16035 10440 16271
rect 10676 16035 10761 16271
rect 10997 16035 11082 16271
rect 11318 16035 11403 16271
rect 11639 16035 11724 16271
rect 11960 16035 12045 16271
rect 12281 16035 12366 16271
rect 12602 16035 12687 16271
rect 12923 16035 13008 16271
rect 13244 16035 13329 16271
rect 13565 16035 13650 16271
rect 13886 16035 13971 16271
rect 14207 16035 14292 16271
rect 14528 16035 14613 16271
rect 14849 16035 15008 16271
rect 8 15935 15008 16035
rect 8 15699 151 15935
rect 387 15699 473 15935
rect 709 15699 795 15935
rect 1031 15699 1117 15935
rect 1353 15699 1439 15935
rect 1675 15699 1761 15935
rect 1997 15699 2083 15935
rect 2319 15699 2405 15935
rect 2641 15699 2727 15935
rect 2963 15699 3049 15935
rect 3285 15699 3371 15935
rect 3607 15699 3693 15935
rect 3929 15699 4015 15935
rect 4251 15699 4337 15935
rect 4573 15699 4659 15935
rect 4895 15699 4981 15935
rect 5217 15699 5303 15935
rect 5539 15699 9477 15935
rect 9713 15699 9798 15935
rect 10034 15699 10119 15935
rect 10355 15699 10440 15935
rect 10676 15699 10761 15935
rect 10997 15699 11082 15935
rect 11318 15699 11403 15935
rect 11639 15699 11724 15935
rect 11960 15699 12045 15935
rect 12281 15699 12366 15935
rect 12602 15699 12687 15935
rect 12923 15699 13008 15935
rect 13244 15699 13329 15935
rect 13565 15699 13650 15935
rect 13886 15699 13971 15935
rect 14207 15699 14292 15935
rect 14528 15699 14613 15935
rect 14849 15699 15008 15935
rect 8 15599 15008 15699
rect 8 15363 151 15599
rect 387 15363 473 15599
rect 709 15363 795 15599
rect 1031 15363 1117 15599
rect 1353 15363 1439 15599
rect 1675 15363 1761 15599
rect 1997 15363 2083 15599
rect 2319 15363 2405 15599
rect 2641 15363 2727 15599
rect 2963 15363 3049 15599
rect 3285 15363 3371 15599
rect 3607 15363 3693 15599
rect 3929 15363 4015 15599
rect 4251 15363 4337 15599
rect 4573 15363 4659 15599
rect 4895 15363 4981 15599
rect 5217 15363 5303 15599
rect 5539 15363 9477 15599
rect 9713 15363 9798 15599
rect 10034 15363 10119 15599
rect 10355 15363 10440 15599
rect 10676 15363 10761 15599
rect 10997 15363 11082 15599
rect 11318 15363 11403 15599
rect 11639 15363 11724 15599
rect 11960 15363 12045 15599
rect 12281 15363 12366 15599
rect 12602 15363 12687 15599
rect 12923 15363 13008 15599
rect 13244 15363 13329 15599
rect 13565 15363 13650 15599
rect 13886 15363 13971 15599
rect 14207 15363 14292 15599
rect 14528 15363 14613 15599
rect 14849 15363 15008 15599
rect 8 15263 15008 15363
rect 8 15027 151 15263
rect 387 15027 473 15263
rect 709 15027 795 15263
rect 1031 15027 1117 15263
rect 1353 15027 1439 15263
rect 1675 15027 1761 15263
rect 1997 15027 2083 15263
rect 2319 15027 2405 15263
rect 2641 15027 2727 15263
rect 2963 15027 3049 15263
rect 3285 15027 3371 15263
rect 3607 15027 3693 15263
rect 3929 15027 4015 15263
rect 4251 15027 4337 15263
rect 4573 15027 4659 15263
rect 4895 15027 4981 15263
rect 5217 15027 5303 15263
rect 5539 15027 9477 15263
rect 9713 15027 9798 15263
rect 10034 15027 10119 15263
rect 10355 15027 10440 15263
rect 10676 15027 10761 15263
rect 10997 15027 11082 15263
rect 11318 15027 11403 15263
rect 11639 15027 11724 15263
rect 11960 15027 12045 15263
rect 12281 15027 12366 15263
rect 12602 15027 12687 15263
rect 12923 15027 13008 15263
rect 13244 15027 13329 15263
rect 13565 15027 13650 15263
rect 13886 15027 13971 15263
rect 14207 15027 14292 15263
rect 14528 15027 14613 15263
rect 14849 15027 15008 15263
rect 8 14927 15008 15027
rect 8 14691 151 14927
rect 387 14691 473 14927
rect 709 14691 795 14927
rect 1031 14691 1117 14927
rect 1353 14691 1439 14927
rect 1675 14691 1761 14927
rect 1997 14691 2083 14927
rect 2319 14691 2405 14927
rect 2641 14691 2727 14927
rect 2963 14691 3049 14927
rect 3285 14691 3371 14927
rect 3607 14691 3693 14927
rect 3929 14691 4015 14927
rect 4251 14691 4337 14927
rect 4573 14691 4659 14927
rect 4895 14691 4981 14927
rect 5217 14691 5303 14927
rect 5539 14691 9477 14927
rect 9713 14691 9798 14927
rect 10034 14691 10119 14927
rect 10355 14691 10440 14927
rect 10676 14691 10761 14927
rect 10997 14691 11082 14927
rect 11318 14691 11403 14927
rect 11639 14691 11724 14927
rect 11960 14691 12045 14927
rect 12281 14691 12366 14927
rect 12602 14691 12687 14927
rect 12923 14691 13008 14927
rect 13244 14691 13329 14927
rect 13565 14691 13650 14927
rect 13886 14691 13971 14927
rect 14207 14691 14292 14927
rect 14528 14691 14613 14927
rect 14849 14691 15008 14927
rect 8 14591 15008 14691
rect 8 14355 151 14591
rect 387 14355 473 14591
rect 709 14355 795 14591
rect 1031 14355 1117 14591
rect 1353 14355 1439 14591
rect 1675 14355 1761 14591
rect 1997 14355 2083 14591
rect 2319 14355 2405 14591
rect 2641 14355 2727 14591
rect 2963 14355 3049 14591
rect 3285 14355 3371 14591
rect 3607 14355 3693 14591
rect 3929 14355 4015 14591
rect 4251 14355 4337 14591
rect 4573 14355 4659 14591
rect 4895 14355 4981 14591
rect 5217 14355 5303 14591
rect 5539 14355 9477 14591
rect 9713 14355 9798 14591
rect 10034 14355 10119 14591
rect 10355 14355 10440 14591
rect 10676 14355 10761 14591
rect 10997 14355 11082 14591
rect 11318 14355 11403 14591
rect 11639 14355 11724 14591
rect 11960 14355 12045 14591
rect 12281 14355 12366 14591
rect 12602 14355 12687 14591
rect 12923 14355 13008 14591
rect 13244 14355 13329 14591
rect 13565 14355 13650 14591
rect 13886 14355 13971 14591
rect 14207 14355 14292 14591
rect 14528 14355 14613 14591
rect 14849 14355 15008 14591
rect 8 14255 15008 14355
rect 8 14019 151 14255
rect 387 14019 473 14255
rect 709 14019 795 14255
rect 1031 14019 1117 14255
rect 1353 14019 1439 14255
rect 1675 14019 1761 14255
rect 1997 14019 2083 14255
rect 2319 14019 2405 14255
rect 2641 14019 2727 14255
rect 2963 14019 3049 14255
rect 3285 14019 3371 14255
rect 3607 14019 3693 14255
rect 3929 14019 4015 14255
rect 4251 14019 4337 14255
rect 4573 14019 4659 14255
rect 4895 14019 4981 14255
rect 5217 14019 5303 14255
rect 5539 14019 9477 14255
rect 9713 14019 9798 14255
rect 10034 14019 10119 14255
rect 10355 14019 10440 14255
rect 10676 14019 10761 14255
rect 10997 14019 11082 14255
rect 11318 14019 11403 14255
rect 11639 14019 11724 14255
rect 11960 14019 12045 14255
rect 12281 14019 12366 14255
rect 12602 14019 12687 14255
rect 12923 14019 13008 14255
rect 13244 14019 13329 14255
rect 13565 14019 13650 14255
rect 13886 14019 13971 14255
rect 14207 14019 14292 14255
rect 14528 14019 14613 14255
rect 14849 14019 15008 14255
rect 8 13994 15008 14019
use sky130_fd_io__pad_esd  sky130_fd_io__pad_esd_0
timestamp 1686671242
transform 1 0 7 0 1 536
box 960 18991 14040 34071
<< labels >>
flabel metal4 s 8 35144 262 39987 3 FreeSans 650 0 0 0 VSSIO
flabel metal4 s 14754 35144 15008 39987 3 FreeSans 650 180 0 0 VSSIO
flabel metal5 s 8 13994 262 18984 3 FreeSans 650 0 0 0 VDDIO
flabel metal4 s 8 13994 262 18987 3 FreeSans 650 0 0 0 VDDIO
flabel metal5 s 14754 13994 15008 18984 3 FreeSans 650 180 0 0 VDDIO
flabel metal4 s 14754 13994 15008 18987 3 FreeSans 650 180 0 0 VDDIO
<< properties >>
string GDS_END 5766170
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 5688624
<< end >>
