magic
tech sky130A
timestamp 1686671242
<< properties >>
string GDS_END 30672382
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30671930
<< end >>
