magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< obsli1 >>
rect 34 2692 2758 2758
rect 34 100 100 2692
rect 260 2466 2532 2532
rect 260 326 326 2466
rect 662 2064 2130 2130
rect 662 728 728 2064
rect 921 921 1871 1871
rect 2064 728 2130 2064
rect 662 662 2130 728
rect 2466 326 2532 2466
rect 260 260 2532 326
rect 2692 100 2758 2692
rect 34 34 2758 100
<< obsm1 >>
rect 38 2696 2754 2754
rect 38 96 96 2696
rect 264 2470 2528 2528
rect 264 322 322 2470
rect 666 2068 2126 2126
rect 666 724 724 2068
rect 935 935 1857 1857
rect 2068 724 2126 2068
rect 666 666 2126 724
rect 2470 322 2528 2470
rect 264 264 2528 322
rect 2696 96 2754 2696
rect 38 38 2754 96
<< properties >>
string FIXED_BBOX 26 26 2766 2766
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9004638
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8927122
<< end >>
