magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 2 21 1839 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 363 47 393 177
rect 447 47 477 177
rect 531 47 561 177
rect 615 47 645 177
rect 699 47 729 177
rect 783 47 813 177
rect 867 47 897 177
rect 951 47 981 177
rect 1139 47 1169 177
rect 1223 47 1253 177
rect 1307 47 1337 177
rect 1391 47 1421 177
rect 1475 47 1505 177
rect 1559 47 1589 177
rect 1643 47 1673 177
rect 1727 47 1757 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 363 297 393 497
rect 447 297 477 497
rect 531 297 561 497
rect 615 297 645 497
rect 699 297 729 497
rect 783 297 813 497
rect 867 297 897 497
rect 951 297 981 497
rect 1139 297 1169 497
rect 1223 297 1253 497
rect 1307 297 1337 497
rect 1391 297 1421 497
rect 1475 297 1505 497
rect 1559 297 1589 497
rect 1643 297 1673 497
rect 1727 297 1757 497
<< ndiff >>
rect 28 163 83 177
rect 28 129 39 163
rect 73 129 83 163
rect 28 95 83 129
rect 28 61 39 95
rect 73 61 83 95
rect 28 47 83 61
rect 113 95 167 177
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 163 249 177
rect 197 129 207 163
rect 241 129 249 163
rect 197 95 249 129
rect 197 61 207 95
rect 241 61 249 95
rect 197 47 249 61
rect 311 95 363 177
rect 311 61 319 95
rect 353 61 363 95
rect 311 47 363 61
rect 393 163 447 177
rect 393 129 403 163
rect 437 129 447 163
rect 393 95 447 129
rect 393 61 403 95
rect 437 61 447 95
rect 393 47 447 61
rect 477 95 531 177
rect 477 61 487 95
rect 521 61 531 95
rect 477 47 531 61
rect 561 163 615 177
rect 561 129 571 163
rect 605 129 615 163
rect 561 95 615 129
rect 561 61 571 95
rect 605 61 615 95
rect 561 47 615 61
rect 645 95 699 177
rect 645 61 655 95
rect 689 61 699 95
rect 645 47 699 61
rect 729 163 783 177
rect 729 129 739 163
rect 773 129 783 163
rect 729 95 783 129
rect 729 61 739 95
rect 773 61 783 95
rect 729 47 783 61
rect 813 95 867 177
rect 813 61 823 95
rect 857 61 867 95
rect 813 47 867 61
rect 897 163 951 177
rect 897 129 907 163
rect 941 129 951 163
rect 897 95 951 129
rect 897 61 907 95
rect 941 61 951 95
rect 897 47 951 61
rect 981 95 1139 177
rect 981 61 991 95
rect 1025 61 1095 95
rect 1129 61 1139 95
rect 981 47 1139 61
rect 1169 163 1223 177
rect 1169 129 1179 163
rect 1213 129 1223 163
rect 1169 95 1223 129
rect 1169 61 1179 95
rect 1213 61 1223 95
rect 1169 47 1223 61
rect 1253 95 1307 177
rect 1253 61 1263 95
rect 1297 61 1307 95
rect 1253 47 1307 61
rect 1337 163 1391 177
rect 1337 129 1347 163
rect 1381 129 1391 163
rect 1337 95 1391 129
rect 1337 61 1347 95
rect 1381 61 1391 95
rect 1337 47 1391 61
rect 1421 95 1475 177
rect 1421 61 1431 95
rect 1465 61 1475 95
rect 1421 47 1475 61
rect 1505 163 1559 177
rect 1505 129 1515 163
rect 1549 129 1559 163
rect 1505 95 1559 129
rect 1505 61 1515 95
rect 1549 61 1559 95
rect 1505 47 1559 61
rect 1589 95 1643 177
rect 1589 61 1599 95
rect 1633 61 1643 95
rect 1589 47 1643 61
rect 1673 163 1727 177
rect 1673 129 1683 163
rect 1717 129 1727 163
rect 1673 95 1727 129
rect 1673 61 1683 95
rect 1717 61 1727 95
rect 1673 47 1727 61
rect 1757 163 1813 177
rect 1757 129 1767 163
rect 1801 129 1813 163
rect 1757 95 1813 129
rect 1757 61 1767 95
rect 1801 61 1813 95
rect 1757 47 1813 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 477 167 497
rect 113 443 123 477
rect 157 443 167 477
rect 113 297 167 443
rect 197 341 253 497
rect 197 307 207 341
rect 241 307 253 341
rect 197 297 253 307
rect 311 477 363 497
rect 311 443 319 477
rect 353 443 363 477
rect 311 297 363 443
rect 393 341 447 497
rect 393 307 403 341
rect 437 307 447 341
rect 393 297 447 307
rect 477 477 531 497
rect 477 443 487 477
rect 521 443 531 477
rect 477 297 531 443
rect 561 341 615 497
rect 561 307 571 341
rect 605 307 615 341
rect 561 297 615 307
rect 645 477 699 497
rect 645 443 655 477
rect 689 443 699 477
rect 645 297 699 443
rect 729 409 783 497
rect 729 375 739 409
rect 773 375 783 409
rect 729 341 783 375
rect 729 307 739 341
rect 773 307 783 341
rect 729 297 783 307
rect 813 477 867 497
rect 813 443 823 477
rect 857 443 867 477
rect 813 409 867 443
rect 813 375 823 409
rect 857 375 867 409
rect 813 297 867 375
rect 897 409 951 497
rect 897 375 907 409
rect 941 375 951 409
rect 897 341 951 375
rect 897 307 907 341
rect 941 307 951 341
rect 897 297 951 307
rect 981 477 1033 497
rect 981 443 991 477
rect 1025 443 1033 477
rect 981 409 1033 443
rect 981 375 991 409
rect 1025 375 1033 409
rect 981 297 1033 375
rect 1087 477 1139 497
rect 1087 443 1095 477
rect 1129 443 1139 477
rect 1087 409 1139 443
rect 1087 375 1095 409
rect 1129 375 1139 409
rect 1087 297 1139 375
rect 1169 409 1223 497
rect 1169 375 1179 409
rect 1213 375 1223 409
rect 1169 341 1223 375
rect 1169 307 1179 341
rect 1213 307 1223 341
rect 1169 297 1223 307
rect 1253 477 1307 497
rect 1253 443 1263 477
rect 1297 443 1307 477
rect 1253 409 1307 443
rect 1253 375 1263 409
rect 1297 375 1307 409
rect 1253 297 1307 375
rect 1337 409 1391 497
rect 1337 375 1347 409
rect 1381 375 1391 409
rect 1337 341 1391 375
rect 1337 307 1347 341
rect 1381 307 1391 341
rect 1337 297 1391 307
rect 1421 477 1475 497
rect 1421 443 1431 477
rect 1465 443 1475 477
rect 1421 409 1475 443
rect 1421 375 1431 409
rect 1465 375 1475 409
rect 1421 341 1475 375
rect 1421 307 1431 341
rect 1465 307 1475 341
rect 1421 297 1475 307
rect 1505 477 1559 497
rect 1505 443 1515 477
rect 1549 443 1559 477
rect 1505 409 1559 443
rect 1505 375 1515 409
rect 1549 375 1559 409
rect 1505 297 1559 375
rect 1589 477 1643 497
rect 1589 443 1599 477
rect 1633 443 1643 477
rect 1589 409 1643 443
rect 1589 375 1599 409
rect 1633 375 1643 409
rect 1589 341 1643 375
rect 1589 307 1599 341
rect 1633 307 1643 341
rect 1589 297 1643 307
rect 1673 477 1727 497
rect 1673 443 1683 477
rect 1717 443 1727 477
rect 1673 409 1727 443
rect 1673 375 1683 409
rect 1717 375 1727 409
rect 1673 297 1727 375
rect 1757 477 1813 497
rect 1757 443 1767 477
rect 1801 443 1813 477
rect 1757 409 1813 443
rect 1757 375 1767 409
rect 1801 375 1813 409
rect 1757 341 1813 375
rect 1757 307 1767 341
rect 1801 307 1813 341
rect 1757 297 1813 307
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 61 157 95
rect 207 129 241 163
rect 207 61 241 95
rect 319 61 353 95
rect 403 129 437 163
rect 403 61 437 95
rect 487 61 521 95
rect 571 129 605 163
rect 571 61 605 95
rect 655 61 689 95
rect 739 129 773 163
rect 739 61 773 95
rect 823 61 857 95
rect 907 129 941 163
rect 907 61 941 95
rect 991 61 1025 95
rect 1095 61 1129 95
rect 1179 129 1213 163
rect 1179 61 1213 95
rect 1263 61 1297 95
rect 1347 129 1381 163
rect 1347 61 1381 95
rect 1431 61 1465 95
rect 1515 129 1549 163
rect 1515 61 1549 95
rect 1599 61 1633 95
rect 1683 129 1717 163
rect 1683 61 1717 95
rect 1767 129 1801 163
rect 1767 61 1801 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 443 157 477
rect 207 307 241 341
rect 319 443 353 477
rect 403 307 437 341
rect 487 443 521 477
rect 571 307 605 341
rect 655 443 689 477
rect 739 375 773 409
rect 739 307 773 341
rect 823 443 857 477
rect 823 375 857 409
rect 907 375 941 409
rect 907 307 941 341
rect 991 443 1025 477
rect 991 375 1025 409
rect 1095 443 1129 477
rect 1095 375 1129 409
rect 1179 375 1213 409
rect 1179 307 1213 341
rect 1263 443 1297 477
rect 1263 375 1297 409
rect 1347 375 1381 409
rect 1347 307 1381 341
rect 1431 443 1465 477
rect 1431 375 1465 409
rect 1431 307 1465 341
rect 1515 443 1549 477
rect 1515 375 1549 409
rect 1599 443 1633 477
rect 1599 375 1633 409
rect 1599 307 1633 341
rect 1683 443 1717 477
rect 1683 375 1717 409
rect 1767 443 1801 477
rect 1767 375 1801 409
rect 1767 307 1801 341
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 363 497 393 523
rect 447 497 477 523
rect 531 497 561 523
rect 615 497 645 523
rect 699 497 729 523
rect 783 497 813 523
rect 867 497 897 523
rect 951 497 981 523
rect 1139 497 1169 523
rect 1223 497 1253 523
rect 1307 497 1337 523
rect 1391 497 1421 523
rect 1475 497 1505 523
rect 1559 497 1589 523
rect 1643 497 1673 523
rect 1727 497 1757 523
rect 83 265 113 297
rect 29 249 113 265
rect 29 215 39 249
rect 73 215 113 249
rect 29 199 113 215
rect 83 177 113 199
rect 167 265 197 297
rect 363 265 393 297
rect 447 265 477 297
rect 531 265 561 297
rect 615 265 645 297
rect 167 249 257 265
rect 167 215 207 249
rect 241 215 257 249
rect 167 199 257 215
rect 363 249 645 265
rect 363 215 383 249
rect 417 215 451 249
rect 485 215 519 249
rect 553 215 645 249
rect 363 199 645 215
rect 167 177 197 199
rect 363 177 393 199
rect 447 177 477 199
rect 531 177 561 199
rect 615 177 645 199
rect 699 265 729 297
rect 783 265 813 297
rect 867 265 897 297
rect 951 265 981 297
rect 699 249 981 265
rect 699 215 727 249
rect 761 215 795 249
rect 829 215 863 249
rect 897 215 931 249
rect 965 215 981 249
rect 699 199 981 215
rect 699 177 729 199
rect 783 177 813 199
rect 867 177 897 199
rect 951 177 981 199
rect 1139 265 1169 297
rect 1223 265 1253 297
rect 1307 265 1337 297
rect 1391 265 1421 297
rect 1139 249 1421 265
rect 1139 215 1167 249
rect 1201 215 1235 249
rect 1269 215 1303 249
rect 1337 215 1371 249
rect 1405 215 1421 249
rect 1139 199 1421 215
rect 1139 177 1169 199
rect 1223 177 1253 199
rect 1307 177 1337 199
rect 1391 177 1421 199
rect 1475 265 1505 297
rect 1559 265 1589 297
rect 1643 265 1673 297
rect 1727 265 1757 297
rect 1475 249 1757 265
rect 1475 215 1503 249
rect 1537 215 1571 249
rect 1605 215 1639 249
rect 1673 215 1707 249
rect 1741 215 1757 249
rect 1475 199 1757 215
rect 1475 177 1505 199
rect 1559 177 1589 199
rect 1643 177 1673 199
rect 1727 177 1757 199
rect 83 21 113 47
rect 167 21 197 47
rect 363 21 393 47
rect 447 21 477 47
rect 531 21 561 47
rect 615 21 645 47
rect 699 21 729 47
rect 783 21 813 47
rect 867 21 897 47
rect 951 21 981 47
rect 1139 21 1169 47
rect 1223 21 1253 47
rect 1307 21 1337 47
rect 1391 21 1421 47
rect 1475 21 1505 47
rect 1559 21 1589 47
rect 1643 21 1673 47
rect 1727 21 1757 47
<< polycont >>
rect 39 215 73 249
rect 207 215 241 249
rect 383 215 417 249
rect 451 215 485 249
rect 519 215 553 249
rect 727 215 761 249
rect 795 215 829 249
rect 863 215 897 249
rect 931 215 965 249
rect 1167 215 1201 249
rect 1235 215 1269 249
rect 1303 215 1337 249
rect 1371 215 1405 249
rect 1503 215 1537 249
rect 1571 215 1605 249
rect 1639 215 1673 249
rect 1707 215 1741 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 17 477 73 493
rect 17 443 39 477
rect 107 477 173 527
rect 107 443 123 477
rect 157 443 173 477
rect 303 477 1039 493
rect 303 443 319 477
rect 353 443 487 477
rect 521 443 655 477
rect 689 459 823 477
rect 689 443 705 459
rect 815 443 823 459
rect 857 459 991 477
rect 857 443 865 459
rect 17 409 73 443
rect 739 409 781 425
rect 17 375 39 409
rect 73 375 705 409
rect 17 341 157 375
rect 17 307 39 341
rect 73 307 157 341
rect 191 307 207 341
rect 241 307 327 341
rect 22 249 89 273
rect 22 215 39 249
rect 73 215 89 249
rect 123 179 157 307
rect 191 249 259 265
rect 191 215 207 249
rect 241 215 259 249
rect 293 249 327 307
rect 368 307 403 341
rect 437 307 571 341
rect 605 307 637 341
rect 368 283 637 307
rect 293 215 383 249
rect 417 215 451 249
rect 485 215 519 249
rect 553 215 569 249
rect 293 181 327 215
rect 603 181 637 283
rect 671 257 705 375
rect 773 375 781 409
rect 739 341 781 375
rect 815 409 865 443
rect 983 443 991 459
rect 1025 443 1039 477
rect 815 375 823 409
rect 857 375 865 409
rect 815 359 865 375
rect 899 409 949 425
rect 899 375 907 409
rect 941 375 949 409
rect 773 325 781 341
rect 899 341 949 375
rect 983 409 1039 443
rect 983 375 991 409
rect 1025 375 1039 409
rect 983 359 1039 375
rect 1076 477 1473 493
rect 1076 443 1095 477
rect 1129 459 1263 477
rect 1129 443 1137 459
rect 1076 409 1137 443
rect 1255 443 1263 459
rect 1297 459 1431 477
rect 1297 443 1305 459
rect 1076 375 1095 409
rect 1129 375 1137 409
rect 1076 359 1137 375
rect 1171 409 1221 425
rect 1171 375 1179 409
rect 1213 375 1221 409
rect 899 325 907 341
rect 773 307 907 325
rect 941 325 949 341
rect 1171 341 1221 375
rect 1255 409 1305 443
rect 1423 443 1431 459
rect 1465 443 1473 477
rect 1255 375 1263 409
rect 1297 375 1305 409
rect 1255 359 1305 375
rect 1339 409 1389 425
rect 1339 375 1347 409
rect 1381 375 1389 409
rect 1171 325 1179 341
rect 941 307 1179 325
rect 1213 325 1221 341
rect 1339 341 1389 375
rect 1339 325 1347 341
rect 1213 307 1347 325
rect 1381 307 1389 341
rect 739 291 1389 307
rect 1423 409 1473 443
rect 1423 375 1431 409
rect 1465 375 1473 409
rect 1423 341 1473 375
rect 1507 477 1557 527
rect 1507 443 1515 477
rect 1549 443 1557 477
rect 1507 409 1557 443
rect 1507 375 1515 409
rect 1549 375 1557 409
rect 1507 359 1557 375
rect 1591 477 1641 493
rect 1591 443 1599 477
rect 1633 443 1641 477
rect 1591 409 1641 443
rect 1591 375 1599 409
rect 1633 375 1641 409
rect 1423 307 1431 341
rect 1465 325 1473 341
rect 1591 341 1641 375
rect 1675 477 1725 527
rect 1675 443 1683 477
rect 1717 443 1725 477
rect 1675 409 1725 443
rect 1675 375 1683 409
rect 1717 375 1725 409
rect 1675 359 1725 375
rect 1759 477 1822 493
rect 1759 443 1767 477
rect 1801 443 1822 477
rect 1759 409 1822 443
rect 1759 375 1767 409
rect 1801 375 1822 409
rect 1591 325 1599 341
rect 1465 307 1599 325
rect 1633 325 1641 341
rect 1759 341 1822 375
rect 1759 325 1767 341
rect 1633 307 1767 325
rect 1801 307 1822 341
rect 1423 291 1822 307
rect 671 249 981 257
rect 671 215 727 249
rect 761 215 795 249
rect 829 215 863 249
rect 897 215 931 249
rect 965 215 981 249
rect 1030 249 1421 257
rect 1030 215 1167 249
rect 1201 215 1235 249
rect 1269 215 1303 249
rect 1337 215 1371 249
rect 1405 215 1421 249
rect 1475 249 1822 257
rect 1475 215 1503 249
rect 1537 215 1571 249
rect 1605 215 1639 249
rect 1673 215 1707 249
rect 1741 215 1822 249
rect 17 163 157 179
rect 17 129 39 163
rect 73 145 157 163
rect 191 163 327 181
rect 73 129 89 145
rect 17 95 89 129
rect 191 129 207 163
rect 241 147 327 163
rect 387 163 1733 181
rect 241 129 257 147
rect 17 61 39 95
rect 73 61 89 95
rect 17 51 89 61
rect 123 95 157 111
rect 123 17 157 61
rect 191 95 257 129
rect 387 129 403 163
rect 437 145 571 163
rect 437 129 453 145
rect 191 61 207 95
rect 241 61 257 95
rect 191 51 257 61
rect 319 95 353 111
rect 319 17 353 61
rect 387 95 453 129
rect 555 129 571 145
rect 605 145 739 163
rect 605 129 621 145
rect 387 61 403 95
rect 437 61 453 95
rect 387 51 453 61
rect 487 95 521 111
rect 487 17 521 61
rect 555 95 621 129
rect 723 129 739 145
rect 773 145 907 163
rect 773 129 789 145
rect 555 61 571 95
rect 605 61 621 95
rect 555 51 621 61
rect 655 95 689 111
rect 655 17 689 61
rect 723 95 789 129
rect 891 129 907 145
rect 941 145 1179 163
rect 941 129 957 145
rect 723 61 739 95
rect 773 61 789 95
rect 723 51 789 61
rect 823 95 857 111
rect 823 17 857 61
rect 891 95 957 129
rect 1163 129 1179 145
rect 1213 145 1347 163
rect 1213 129 1229 145
rect 891 61 907 95
rect 941 61 957 95
rect 891 51 957 61
rect 991 95 1129 111
rect 1025 61 1095 95
rect 991 17 1129 61
rect 1163 95 1229 129
rect 1331 129 1347 145
rect 1381 145 1515 163
rect 1381 129 1397 145
rect 1163 61 1179 95
rect 1213 61 1229 95
rect 1163 51 1229 61
rect 1263 95 1297 111
rect 1263 17 1297 61
rect 1331 95 1397 129
rect 1499 129 1515 145
rect 1549 145 1683 163
rect 1549 129 1565 145
rect 1331 61 1347 95
rect 1381 61 1397 95
rect 1331 51 1397 61
rect 1431 95 1465 111
rect 1431 17 1465 61
rect 1499 95 1565 129
rect 1667 129 1683 145
rect 1717 129 1733 163
rect 1499 61 1515 95
rect 1549 61 1565 95
rect 1499 51 1565 61
rect 1599 95 1633 111
rect 1599 17 1633 61
rect 1667 95 1733 129
rect 1667 61 1683 95
rect 1717 61 1733 95
rect 1667 51 1733 61
rect 1767 163 1822 181
rect 1801 129 1822 163
rect 1767 95 1822 129
rect 1801 61 1822 95
rect 1767 17 1822 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel locali s 214 221 248 255 0 FreeSans 400 180 0 0 D_N
port 4 nsew signal input
flabel locali s 580 289 614 323 0 FreeSans 400 180 0 0 Y
port 9 nsew signal output
flabel locali s 1592 221 1626 255 0 FreeSans 400 180 0 0 A
port 1 nsew signal input
flabel locali s 1224 221 1258 255 0 FreeSans 400 180 0 0 B
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel mvpsubdiff s 38 61 38 61 0 FreeSans 240 0 0 0 k
rlabel comment s 0 0 0 0 4 nor4bb_4
rlabel metal1 s 0 -48 1840 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1840 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1840 544
string GDS_END 1210492
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1196968
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 9.200 0.000 
<< end >>
