magic
tech sky130A
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_0
timestamp 1686671242
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 48783660
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48782866
<< end >>
