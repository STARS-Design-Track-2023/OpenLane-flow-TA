magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 314 582
<< pwell >>
rect 1 21 271 203
rect 30 -17 64 21
<< locali >>
rect 19 333 85 490
rect 19 299 155 333
rect 17 215 87 265
rect 121 179 155 299
rect 189 215 259 265
rect 103 51 169 179
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 191 299 257 527
rect 21 17 69 179
rect 203 17 257 179
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
rlabel locali s 189 215 259 265 6 A
port 1 nsew signal input
rlabel locali s 17 215 87 265 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 276 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 271 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 314 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 276 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 103 51 169 179 6 Y
port 7 nsew signal output
rlabel locali s 121 179 155 299 6 Y
port 7 nsew signal output
rlabel locali s 19 299 155 333 6 Y
port 7 nsew signal output
rlabel locali s 19 333 85 490 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 276 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1962442
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1958836
<< end >>
