magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -36 679 1268 1471
<< pwell >>
rect 1096 25 1198 159
<< psubdiff >>
rect 1122 109 1172 133
rect 1122 75 1130 109
rect 1164 75 1172 109
rect 1122 51 1172 75
<< nsubdiff >>
rect 1122 1339 1172 1363
rect 1122 1305 1130 1339
rect 1164 1305 1172 1339
rect 1122 1281 1172 1305
<< psubdiffcont >>
rect 1130 75 1164 109
<< nsubdiffcont >>
rect 1130 1305 1164 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 1232 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1130 1339 1164 1397
rect 1130 1289 1164 1305
rect 64 724 98 740
rect 64 674 98 690
rect 596 724 630 1096
rect 596 690 647 724
rect 596 318 630 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1130 109 1164 125
rect 1130 17 1164 75
rect 0 -17 1232 17
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_16  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_16_0
timestamp 1686671242
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_28  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_28_0
timestamp 1686671242
transform 1 0 1122 0 1 1281
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_29  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_29_0
timestamp 1686671242
transform 1 0 1122 0 1 51
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_nmos_m9_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_8x1024_8_nmos_m9_w2_000_sli_dli_da_p_0
timestamp 1686671242
transform 1 0 54 0 1 51
box -26 -26 1040 456
use sky130_sram_1kbyte_1rw1r_8x1024_8_pmos_m9_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_8x1024_8_pmos_m9_w2_000_sli_dli_da_p_0
timestamp 1686671242
transform 1 0 54 0 1 963
box -59 -56 1073 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 630 707 630 707 4 Z
rlabel locali s 616 0 616 0 4 gnd
rlabel locali s 616 1414 616 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1232 1414
string GDS_END 85032
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 82650
<< end >>
