magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 459 203
rect 30 -17 64 21
<< locali >>
rect 375 333 442 489
rect 214 289 291 333
rect 17 199 73 265
rect 122 67 211 255
rect 254 199 291 289
rect 325 299 442 333
rect 325 165 359 299
rect 393 199 443 265
rect 276 143 359 165
rect 276 59 357 143
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 18 299 84 527
rect 118 401 153 483
rect 187 435 253 527
rect 294 401 339 483
rect 118 367 339 401
rect 18 17 86 163
rect 391 17 443 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 254 199 291 289 6 A1
port 1 nsew signal input
rlabel locali s 214 289 291 333 6 A1
port 1 nsew signal input
rlabel locali s 122 67 211 255 6 A2
port 2 nsew signal input
rlabel locali s 17 199 73 265 6 A3
port 3 nsew signal input
rlabel locali s 393 199 443 265 6 B1
port 4 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 459 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 276 59 357 143 6 Y
port 9 nsew signal output
rlabel locali s 276 143 359 165 6 Y
port 9 nsew signal output
rlabel locali s 325 165 359 299 6 Y
port 9 nsew signal output
rlabel locali s 325 299 442 333 6 Y
port 9 nsew signal output
rlabel locali s 375 333 442 489 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4142840
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4137594
<< end >>
