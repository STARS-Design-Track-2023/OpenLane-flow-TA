magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1555 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 419 47 449 177
rect 503 47 533 177
rect 587 47 617 177
rect 671 47 701 177
rect 859 47 889 177
rect 943 47 973 177
rect 1027 47 1057 177
rect 1111 47 1141 177
rect 1195 47 1225 177
rect 1279 47 1309 177
rect 1363 47 1393 177
rect 1447 47 1477 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 419 297 449 497
rect 503 297 533 497
rect 587 297 617 497
rect 671 297 701 497
rect 859 297 889 497
rect 943 297 973 497
rect 1027 297 1057 497
rect 1111 297 1141 497
rect 1195 297 1225 497
rect 1279 297 1309 497
rect 1363 297 1393 497
rect 1447 297 1477 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 95 335 129
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 95 419 177
rect 365 61 375 95
rect 409 61 419 95
rect 365 47 419 61
rect 449 163 503 177
rect 449 129 459 163
rect 493 129 503 163
rect 449 95 503 129
rect 449 61 459 95
rect 493 61 503 95
rect 449 47 503 61
rect 533 95 587 177
rect 533 61 543 95
rect 577 61 587 95
rect 533 47 587 61
rect 617 163 671 177
rect 617 129 627 163
rect 661 129 671 163
rect 617 95 671 129
rect 617 61 627 95
rect 661 61 671 95
rect 617 47 671 61
rect 701 95 859 177
rect 701 61 711 95
rect 745 61 815 95
rect 849 61 859 95
rect 701 47 859 61
rect 889 163 943 177
rect 889 129 899 163
rect 933 129 943 163
rect 889 95 943 129
rect 889 61 899 95
rect 933 61 943 95
rect 889 47 943 61
rect 973 95 1027 177
rect 973 61 983 95
rect 1017 61 1027 95
rect 973 47 1027 61
rect 1057 163 1111 177
rect 1057 129 1067 163
rect 1101 129 1111 163
rect 1057 95 1111 129
rect 1057 61 1067 95
rect 1101 61 1111 95
rect 1057 47 1111 61
rect 1141 95 1195 177
rect 1141 61 1151 95
rect 1185 61 1195 95
rect 1141 47 1195 61
rect 1225 163 1279 177
rect 1225 129 1235 163
rect 1269 129 1279 163
rect 1225 95 1279 129
rect 1225 61 1235 95
rect 1269 61 1279 95
rect 1225 47 1279 61
rect 1309 95 1363 177
rect 1309 61 1319 95
rect 1353 61 1363 95
rect 1309 47 1363 61
rect 1393 163 1447 177
rect 1393 129 1403 163
rect 1437 129 1447 163
rect 1393 95 1447 129
rect 1393 61 1403 95
rect 1437 61 1447 95
rect 1393 47 1447 61
rect 1477 95 1529 177
rect 1477 61 1487 95
rect 1521 61 1529 95
rect 1477 47 1529 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 477 167 497
rect 113 443 123 477
rect 157 443 167 477
rect 113 409 167 443
rect 113 375 123 409
rect 157 375 167 409
rect 113 297 167 375
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 341 251 375
rect 197 307 207 341
rect 241 307 251 341
rect 197 297 251 307
rect 281 477 335 497
rect 281 443 291 477
rect 325 443 335 477
rect 281 409 335 443
rect 281 375 291 409
rect 325 375 335 409
rect 281 297 335 375
rect 365 477 419 497
rect 365 443 375 477
rect 409 443 419 477
rect 365 409 419 443
rect 365 375 375 409
rect 409 375 419 409
rect 365 341 419 375
rect 365 307 375 341
rect 409 307 419 341
rect 365 297 419 307
rect 449 409 503 497
rect 449 375 459 409
rect 493 375 503 409
rect 449 341 503 375
rect 449 307 459 341
rect 493 307 503 341
rect 449 297 503 307
rect 533 477 587 497
rect 533 443 543 477
rect 577 443 587 477
rect 533 409 587 443
rect 533 375 543 409
rect 577 375 587 409
rect 533 297 587 375
rect 617 409 671 497
rect 617 375 627 409
rect 661 375 671 409
rect 617 341 671 375
rect 617 307 627 341
rect 661 307 671 341
rect 617 297 671 307
rect 701 477 753 497
rect 701 443 711 477
rect 745 443 753 477
rect 701 409 753 443
rect 701 375 711 409
rect 745 375 753 409
rect 701 297 753 375
rect 807 477 859 497
rect 807 443 815 477
rect 849 443 859 477
rect 807 409 859 443
rect 807 375 815 409
rect 849 375 859 409
rect 807 297 859 375
rect 889 409 943 497
rect 889 375 899 409
rect 933 375 943 409
rect 889 341 943 375
rect 889 307 899 341
rect 933 307 943 341
rect 889 297 943 307
rect 973 477 1027 497
rect 973 443 983 477
rect 1017 443 1027 477
rect 973 409 1027 443
rect 973 375 983 409
rect 1017 375 1027 409
rect 973 297 1027 375
rect 1057 409 1111 497
rect 1057 375 1067 409
rect 1101 375 1111 409
rect 1057 341 1111 375
rect 1057 307 1067 341
rect 1101 307 1111 341
rect 1057 297 1111 307
rect 1141 477 1195 497
rect 1141 443 1151 477
rect 1185 443 1195 477
rect 1141 409 1195 443
rect 1141 375 1151 409
rect 1185 375 1195 409
rect 1141 297 1195 375
rect 1225 409 1279 497
rect 1225 375 1235 409
rect 1269 375 1279 409
rect 1225 341 1279 375
rect 1225 307 1235 341
rect 1269 307 1279 341
rect 1225 297 1279 307
rect 1309 477 1363 497
rect 1309 443 1319 477
rect 1353 443 1363 477
rect 1309 409 1363 443
rect 1309 375 1319 409
rect 1353 375 1363 409
rect 1309 297 1363 375
rect 1393 409 1447 497
rect 1393 375 1403 409
rect 1437 375 1447 409
rect 1393 341 1447 375
rect 1393 307 1403 341
rect 1437 307 1447 341
rect 1393 297 1447 307
rect 1477 477 1529 497
rect 1477 443 1487 477
rect 1521 443 1529 477
rect 1477 409 1529 443
rect 1477 375 1487 409
rect 1521 375 1529 409
rect 1477 297 1529 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 61 241 95
rect 291 129 325 163
rect 291 61 325 95
rect 375 61 409 95
rect 459 129 493 163
rect 459 61 493 95
rect 543 61 577 95
rect 627 129 661 163
rect 627 61 661 95
rect 711 61 745 95
rect 815 61 849 95
rect 899 129 933 163
rect 899 61 933 95
rect 983 61 1017 95
rect 1067 129 1101 163
rect 1067 61 1101 95
rect 1151 61 1185 95
rect 1235 129 1269 163
rect 1235 61 1269 95
rect 1319 61 1353 95
rect 1403 129 1437 163
rect 1403 61 1437 95
rect 1487 61 1521 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 443 157 477
rect 123 375 157 409
rect 207 443 241 477
rect 207 375 241 409
rect 207 307 241 341
rect 291 443 325 477
rect 291 375 325 409
rect 375 443 409 477
rect 375 375 409 409
rect 375 307 409 341
rect 459 375 493 409
rect 459 307 493 341
rect 543 443 577 477
rect 543 375 577 409
rect 627 375 661 409
rect 627 307 661 341
rect 711 443 745 477
rect 711 375 745 409
rect 815 443 849 477
rect 815 375 849 409
rect 899 375 933 409
rect 899 307 933 341
rect 983 443 1017 477
rect 983 375 1017 409
rect 1067 375 1101 409
rect 1067 307 1101 341
rect 1151 443 1185 477
rect 1151 375 1185 409
rect 1235 375 1269 409
rect 1235 307 1269 341
rect 1319 443 1353 477
rect 1319 375 1353 409
rect 1403 375 1437 409
rect 1403 307 1437 341
rect 1487 443 1521 477
rect 1487 375 1521 409
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 419 497 449 523
rect 503 497 533 523
rect 587 497 617 523
rect 671 497 701 523
rect 859 497 889 523
rect 943 497 973 523
rect 1027 497 1057 523
rect 1111 497 1141 523
rect 1195 497 1225 523
rect 1279 497 1309 523
rect 1363 497 1393 523
rect 1447 497 1477 523
rect 83 265 113 297
rect 167 265 197 297
rect 251 265 281 297
rect 335 265 365 297
rect 83 249 365 265
rect 83 215 99 249
rect 133 215 167 249
rect 201 215 235 249
rect 269 215 303 249
rect 337 215 365 249
rect 83 199 365 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 177 281 199
rect 335 177 365 199
rect 419 265 449 297
rect 503 265 533 297
rect 587 265 617 297
rect 671 265 701 297
rect 419 249 701 265
rect 419 215 435 249
rect 469 215 503 249
rect 537 215 571 249
rect 605 215 639 249
rect 673 215 701 249
rect 419 199 701 215
rect 419 177 449 199
rect 503 177 533 199
rect 587 177 617 199
rect 671 177 701 199
rect 859 265 889 297
rect 943 265 973 297
rect 1027 265 1057 297
rect 1111 265 1141 297
rect 859 249 1141 265
rect 859 215 875 249
rect 909 215 943 249
rect 977 215 1011 249
rect 1045 215 1079 249
rect 1113 215 1141 249
rect 859 199 1141 215
rect 859 177 889 199
rect 943 177 973 199
rect 1027 177 1057 199
rect 1111 177 1141 199
rect 1195 265 1225 297
rect 1279 265 1309 297
rect 1363 265 1393 297
rect 1447 265 1477 297
rect 1195 249 1477 265
rect 1195 215 1205 249
rect 1239 215 1273 249
rect 1307 215 1341 249
rect 1375 215 1409 249
rect 1443 215 1477 249
rect 1195 199 1477 215
rect 1195 177 1225 199
rect 1279 177 1309 199
rect 1363 177 1393 199
rect 1447 177 1477 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 419 21 449 47
rect 503 21 533 47
rect 587 21 617 47
rect 671 21 701 47
rect 859 21 889 47
rect 943 21 973 47
rect 1027 21 1057 47
rect 1111 21 1141 47
rect 1195 21 1225 47
rect 1279 21 1309 47
rect 1363 21 1393 47
rect 1447 21 1477 47
<< polycont >>
rect 99 215 133 249
rect 167 215 201 249
rect 235 215 269 249
rect 303 215 337 249
rect 435 215 469 249
rect 503 215 537 249
rect 571 215 605 249
rect 639 215 673 249
rect 875 215 909 249
rect 943 215 977 249
rect 1011 215 1045 249
rect 1079 215 1113 249
rect 1205 215 1239 249
rect 1273 215 1307 249
rect 1341 215 1375 249
rect 1409 215 1443 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 18 477 81 493
rect 18 443 39 477
rect 73 443 81 477
rect 18 409 81 443
rect 18 375 39 409
rect 73 375 81 409
rect 18 341 81 375
rect 115 477 165 527
rect 115 443 123 477
rect 157 443 165 477
rect 115 409 165 443
rect 115 375 123 409
rect 157 375 165 409
rect 115 359 165 375
rect 199 477 249 493
rect 199 443 207 477
rect 241 443 249 477
rect 199 409 249 443
rect 199 375 207 409
rect 241 375 249 409
rect 18 307 39 341
rect 73 325 81 341
rect 199 341 249 375
rect 283 477 333 527
rect 283 443 291 477
rect 325 443 333 477
rect 283 409 333 443
rect 283 375 291 409
rect 325 375 333 409
rect 283 359 333 375
rect 367 477 764 493
rect 367 443 375 477
rect 409 459 543 477
rect 409 443 417 459
rect 367 409 417 443
rect 535 443 543 459
rect 577 459 711 477
rect 577 443 585 459
rect 367 375 375 409
rect 409 375 417 409
rect 199 325 207 341
rect 73 307 207 325
rect 241 325 249 341
rect 367 341 417 375
rect 367 325 375 341
rect 241 307 375 325
rect 409 307 417 341
rect 18 291 417 307
rect 451 409 501 425
rect 451 375 459 409
rect 493 375 501 409
rect 451 341 501 375
rect 535 409 585 443
rect 703 443 711 459
rect 745 443 764 477
rect 535 375 543 409
rect 577 375 585 409
rect 535 359 585 375
rect 619 409 669 425
rect 619 375 627 409
rect 661 375 669 409
rect 451 307 459 341
rect 493 325 501 341
rect 619 341 669 375
rect 703 409 764 443
rect 703 375 711 409
rect 745 375 764 409
rect 703 359 764 375
rect 801 477 1529 493
rect 801 443 815 477
rect 849 459 983 477
rect 849 443 857 459
rect 801 409 857 443
rect 975 443 983 459
rect 1017 459 1151 477
rect 1017 443 1025 459
rect 801 375 815 409
rect 849 375 857 409
rect 801 359 857 375
rect 891 409 941 425
rect 891 375 899 409
rect 933 375 941 409
rect 619 325 627 341
rect 493 307 627 325
rect 661 325 669 341
rect 891 341 941 375
rect 975 409 1025 443
rect 1143 443 1151 459
rect 1185 459 1319 477
rect 1185 443 1193 459
rect 975 375 983 409
rect 1017 375 1025 409
rect 975 359 1025 375
rect 1059 409 1109 425
rect 1059 375 1067 409
rect 1101 375 1109 409
rect 891 325 899 341
rect 661 307 899 325
rect 933 325 941 341
rect 1059 341 1109 375
rect 1143 409 1193 443
rect 1311 443 1319 459
rect 1353 459 1487 477
rect 1353 443 1361 459
rect 1143 375 1151 409
rect 1185 375 1193 409
rect 1143 359 1193 375
rect 1227 409 1277 425
rect 1227 375 1235 409
rect 1269 375 1277 409
rect 1059 325 1067 341
rect 933 307 1067 325
rect 1101 307 1109 341
rect 451 291 1109 307
rect 1227 341 1277 375
rect 1311 409 1361 443
rect 1479 443 1487 459
rect 1521 443 1529 477
rect 1311 375 1319 409
rect 1353 375 1361 409
rect 1311 359 1361 375
rect 1395 409 1445 425
rect 1395 375 1403 409
rect 1437 375 1445 409
rect 1227 307 1235 341
rect 1269 325 1277 341
rect 1395 341 1445 375
rect 1479 409 1529 443
rect 1479 375 1487 409
rect 1521 375 1529 409
rect 1479 359 1529 375
rect 1395 325 1403 341
rect 1269 307 1403 325
rect 1437 325 1445 341
rect 1437 307 1547 325
rect 1227 291 1547 307
rect 36 249 365 257
rect 36 215 99 249
rect 133 215 167 249
rect 201 215 235 249
rect 269 215 303 249
rect 337 215 365 249
rect 419 249 814 257
rect 419 215 435 249
rect 469 215 503 249
rect 537 215 571 249
rect 605 215 639 249
rect 673 215 814 249
rect 859 249 1141 257
rect 859 215 875 249
rect 909 215 943 249
rect 977 215 1011 249
rect 1045 215 1079 249
rect 1113 215 1141 249
rect 1175 249 1459 257
rect 1175 215 1205 249
rect 1239 215 1273 249
rect 1307 215 1341 249
rect 1375 215 1409 249
rect 1443 215 1459 249
rect 1493 181 1547 291
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 1547 181
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 107 95 173 129
rect 275 129 291 145
rect 325 145 459 163
rect 325 129 341 145
rect 107 61 123 95
rect 157 61 173 95
rect 107 51 173 61
rect 207 95 241 111
rect 207 17 241 61
rect 275 95 341 129
rect 443 129 459 145
rect 493 145 627 163
rect 493 129 509 145
rect 275 61 291 95
rect 325 61 341 95
rect 275 51 341 61
rect 375 95 409 111
rect 375 17 409 61
rect 443 95 509 129
rect 611 129 627 145
rect 661 145 899 163
rect 661 129 677 145
rect 443 61 459 95
rect 493 61 509 95
rect 443 51 509 61
rect 543 95 577 111
rect 543 17 577 61
rect 611 95 677 129
rect 883 129 899 145
rect 933 145 1067 163
rect 933 129 949 145
rect 611 61 627 95
rect 661 61 677 95
rect 611 51 677 61
rect 711 95 849 111
rect 745 61 815 95
rect 711 17 849 61
rect 883 95 949 129
rect 1051 129 1067 145
rect 1101 145 1235 163
rect 1101 129 1117 145
rect 883 61 899 95
rect 933 61 949 95
rect 883 51 949 61
rect 983 95 1017 111
rect 983 17 1017 61
rect 1051 95 1117 129
rect 1219 129 1235 145
rect 1269 145 1403 163
rect 1269 129 1285 145
rect 1051 61 1067 95
rect 1101 61 1117 95
rect 1051 51 1117 61
rect 1151 95 1185 111
rect 1151 17 1185 61
rect 1219 95 1285 129
rect 1387 129 1403 145
rect 1437 145 1547 163
rect 1437 129 1453 145
rect 1219 61 1235 95
rect 1269 61 1285 95
rect 1219 51 1285 61
rect 1319 95 1353 111
rect 1319 17 1353 61
rect 1387 95 1453 129
rect 1387 61 1403 95
rect 1437 61 1453 95
rect 1387 51 1453 61
rect 1487 95 1521 111
rect 1487 17 1521 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 214 221 248 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 950 221 984 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 1502 153 1536 187 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 1318 221 1352 255 0 FreeSans 400 0 0 0 D
port 4 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 766 221 800 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor4_4
rlabel metal1 s 0 -48 1564 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 1152972
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1140654
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 7.820 0.000 
<< end >>
