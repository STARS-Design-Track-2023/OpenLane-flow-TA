magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< locali >>
rect 217 752 255 786
rect 289 752 327 786
rect 361 752 399 786
rect 433 752 471 786
rect 505 752 543 786
rect 577 752 615 786
rect 649 752 687 786
rect 721 752 759 786
rect 48 672 82 674
rect 48 600 82 638
rect 48 528 82 566
rect 48 456 82 494
rect 48 384 82 422
rect 48 312 82 350
rect 48 240 82 278
rect 48 168 82 206
rect 48 132 82 134
rect 894 672 928 674
rect 894 600 928 638
rect 894 528 928 566
rect 894 456 928 494
rect 894 384 928 422
rect 894 312 928 350
rect 894 240 928 278
rect 894 168 928 206
rect 894 132 928 134
rect 217 20 255 54
rect 289 20 327 54
rect 361 20 399 54
rect 433 20 471 54
rect 505 20 543 54
rect 577 20 615 54
rect 649 20 687 54
rect 721 20 759 54
<< viali >>
rect 183 752 217 786
rect 255 752 289 786
rect 327 752 361 786
rect 399 752 433 786
rect 471 752 505 786
rect 543 752 577 786
rect 615 752 649 786
rect 687 752 721 786
rect 759 752 793 786
rect 48 638 82 672
rect 48 566 82 600
rect 48 494 82 528
rect 48 422 82 456
rect 48 350 82 384
rect 48 278 82 312
rect 48 206 82 240
rect 48 134 82 168
rect 894 638 928 672
rect 894 566 928 600
rect 894 494 928 528
rect 894 422 928 456
rect 894 350 928 384
rect 894 278 928 312
rect 894 206 928 240
rect 894 134 928 168
rect 183 20 217 54
rect 255 20 289 54
rect 327 20 361 54
rect 399 20 433 54
rect 471 20 505 54
rect 543 20 577 54
rect 615 20 649 54
rect 687 20 721 54
rect 759 20 793 54
<< obsli1 >>
rect 159 98 193 708
rect 315 98 349 708
rect 471 98 505 708
rect 627 98 661 708
rect 783 98 817 708
<< metal1 >>
rect 171 786 805 806
rect 171 752 183 786
rect 217 752 255 786
rect 289 752 327 786
rect 361 752 399 786
rect 433 752 471 786
rect 505 752 543 786
rect 577 752 615 786
rect 649 752 687 786
rect 721 752 759 786
rect 793 752 805 786
rect 171 740 805 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 882 672 940 684
rect 882 638 894 672
rect 928 638 940 672
rect 882 600 940 638
rect 882 566 894 600
rect 928 566 940 600
rect 882 528 940 566
rect 882 494 894 528
rect 928 494 940 528
rect 882 456 940 494
rect 882 422 894 456
rect 928 422 940 456
rect 882 384 940 422
rect 882 350 894 384
rect 928 350 940 384
rect 882 312 940 350
rect 882 278 894 312
rect 928 278 940 312
rect 882 240 940 278
rect 882 206 894 240
rect 928 206 940 240
rect 882 168 940 206
rect 882 134 894 168
rect 928 134 940 168
rect 882 122 940 134
rect 171 54 805 66
rect 171 20 183 54
rect 217 20 255 54
rect 289 20 327 54
rect 361 20 399 54
rect 433 20 471 54
rect 505 20 543 54
rect 577 20 615 54
rect 649 20 687 54
rect 721 20 759 54
rect 793 20 805 54
rect 171 0 805 20
<< obsm1 >>
rect 150 122 202 684
rect 306 122 358 684
rect 462 122 514 684
rect 618 122 670 684
rect 774 122 826 684
<< metal2 >>
rect 10 428 966 684
rect 10 122 966 378
<< labels >>
rlabel viali s 894 638 928 672 6 BULK
port 1 nsew
rlabel viali s 894 566 928 600 6 BULK
port 1 nsew
rlabel viali s 894 494 928 528 6 BULK
port 1 nsew
rlabel viali s 894 422 928 456 6 BULK
port 1 nsew
rlabel viali s 894 350 928 384 6 BULK
port 1 nsew
rlabel viali s 894 278 928 312 6 BULK
port 1 nsew
rlabel viali s 894 206 928 240 6 BULK
port 1 nsew
rlabel viali s 894 134 928 168 6 BULK
port 1 nsew
rlabel viali s 48 638 82 672 6 BULK
port 1 nsew
rlabel viali s 48 566 82 600 6 BULK
port 1 nsew
rlabel viali s 48 494 82 528 6 BULK
port 1 nsew
rlabel viali s 48 422 82 456 6 BULK
port 1 nsew
rlabel viali s 48 350 82 384 6 BULK
port 1 nsew
rlabel viali s 48 278 82 312 6 BULK
port 1 nsew
rlabel viali s 48 206 82 240 6 BULK
port 1 nsew
rlabel viali s 48 134 82 168 6 BULK
port 1 nsew
rlabel locali s 894 132 928 674 6 BULK
port 1 nsew
rlabel locali s 48 132 82 674 6 BULK
port 1 nsew
rlabel metal1 s 882 122 940 684 6 BULK
port 1 nsew
rlabel metal1 s 36 122 94 684 6 BULK
port 1 nsew
rlabel metal2 s 10 428 966 684 6 DRAIN
port 2 nsew
rlabel viali s 759 752 793 786 6 GATE
port 3 nsew
rlabel viali s 759 20 793 54 6 GATE
port 3 nsew
rlabel viali s 687 752 721 786 6 GATE
port 3 nsew
rlabel viali s 687 20 721 54 6 GATE
port 3 nsew
rlabel viali s 615 752 649 786 6 GATE
port 3 nsew
rlabel viali s 615 20 649 54 6 GATE
port 3 nsew
rlabel viali s 543 752 577 786 6 GATE
port 3 nsew
rlabel viali s 543 20 577 54 6 GATE
port 3 nsew
rlabel viali s 471 752 505 786 6 GATE
port 3 nsew
rlabel viali s 471 20 505 54 6 GATE
port 3 nsew
rlabel viali s 399 752 433 786 6 GATE
port 3 nsew
rlabel viali s 399 20 433 54 6 GATE
port 3 nsew
rlabel viali s 327 752 361 786 6 GATE
port 3 nsew
rlabel viali s 327 20 361 54 6 GATE
port 3 nsew
rlabel viali s 255 752 289 786 6 GATE
port 3 nsew
rlabel viali s 255 20 289 54 6 GATE
port 3 nsew
rlabel viali s 183 752 217 786 6 GATE
port 3 nsew
rlabel viali s 183 20 217 54 6 GATE
port 3 nsew
rlabel locali s 183 752 793 786 6 GATE
port 3 nsew
rlabel locali s 183 20 793 54 6 GATE
port 3 nsew
rlabel metal1 s 171 740 805 806 6 GATE
port 3 nsew
rlabel metal1 s 171 0 805 66 6 GATE
port 3 nsew
rlabel metal2 s 10 122 966 378 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 976 806
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9963674
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9947658
<< end >>
