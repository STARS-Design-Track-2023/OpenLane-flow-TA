magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -66 377 738 897
<< pwell >>
rect 50 43 668 283
rect -26 -43 698 43
<< locali >>
rect 240 356 274 751
rect 25 344 274 356
rect 409 355 555 424
rect 25 310 278 344
rect 244 99 278 310
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 18 735 204 751
rect 18 701 22 735
rect 56 701 94 735
rect 128 701 166 735
rect 200 701 204 735
rect 18 435 204 701
rect 310 735 560 751
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 310 460 560 701
rect 18 113 208 265
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 208 113
rect 314 319 373 351
rect 596 319 650 601
rect 314 285 650 319
rect 314 113 564 249
rect 600 165 650 285
rect 18 73 208 79
rect 348 79 386 113
rect 420 79 458 113
rect 492 79 530 113
rect 314 73 564 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 22 701 56 735
rect 94 701 128 735
rect 166 701 200 735
rect 310 701 344 735
rect 382 701 416 735
rect 454 701 488 735
rect 526 701 560 735
rect 24 79 58 113
rect 96 79 130 113
rect 168 79 202 113
rect 314 79 348 113
rect 386 79 420 113
rect 458 79 492 113
rect 530 79 564 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 831 672 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 0 791 672 797
rect 0 735 672 763
rect 0 701 22 735
rect 56 701 94 735
rect 128 701 166 735
rect 200 701 310 735
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 560 701 672 735
rect 0 689 672 701
rect 0 113 672 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 314 113
rect 348 79 386 113
rect 420 79 458 113
rect 492 79 530 113
rect 564 79 672 113
rect 0 51 672 79
rect 0 17 672 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -23 672 -17
<< labels >>
rlabel locali s 409 355 555 424 6 A
port 1 nsew signal input
rlabel metal1 s 0 51 672 125 6 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 -23 672 23 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s -26 -43 698 43 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 50 43 668 283 6 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 791 672 837 6 VPB
port 4 nsew power bidirectional
rlabel nwell s -66 377 738 897 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 689 672 763 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 244 99 278 310 6 X
port 6 nsew signal output
rlabel locali s 25 310 278 344 6 X
port 6 nsew signal output
rlabel locali s 25 344 274 356 6 X
port 6 nsew signal output
rlabel locali s 240 356 274 751 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 672 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 829860
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 821298
<< end >>
