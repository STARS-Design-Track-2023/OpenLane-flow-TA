magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 2430 582
<< pwell >>
rect 1 21 2391 203
rect 30 -17 64 21
<< locali >>
rect 1047 323 1113 493
rect 1215 323 1281 493
rect 1383 323 1449 493
rect 1551 323 1617 493
rect 1719 323 1785 493
rect 1887 323 1953 493
rect 2055 323 2121 493
rect 2223 323 2289 493
rect 1047 289 2375 323
rect 22 215 88 255
rect 2324 181 2375 289
rect 1047 147 2375 181
rect 1047 52 1113 147
rect 1047 51 1097 52
rect 1215 52 1281 147
rect 1231 51 1265 52
rect 1383 52 1449 147
rect 1399 51 1433 52
rect 1551 52 1617 147
rect 1719 52 1785 147
rect 1887 52 1953 147
rect 2055 52 2121 147
rect 2223 52 2289 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 35 289 69 527
rect 103 289 169 493
rect 207 323 273 493
rect 307 357 341 527
rect 375 323 441 493
rect 475 357 509 527
rect 543 323 609 493
rect 643 367 677 527
rect 711 323 777 493
rect 811 367 845 527
rect 879 323 945 493
rect 979 367 1013 527
rect 1147 367 1181 527
rect 1315 367 1349 527
rect 1483 367 1517 527
rect 1651 367 1685 527
rect 1819 367 1853 527
rect 1987 367 2021 527
rect 2155 367 2189 527
rect 2323 367 2357 527
rect 207 289 509 323
rect 543 289 1013 323
rect 122 255 169 289
rect 475 255 509 289
rect 978 255 1013 289
rect 122 215 441 255
rect 475 215 937 255
rect 978 215 2290 255
rect 122 181 169 215
rect 475 181 509 215
rect 978 181 1013 215
rect 35 17 69 181
rect 103 52 169 181
rect 207 147 509 181
rect 543 147 1013 181
rect 207 52 273 147
rect 307 17 341 113
rect 375 52 441 147
rect 475 17 509 113
rect 543 52 609 147
rect 643 17 677 113
rect 711 52 777 147
rect 811 17 845 113
rect 879 52 945 147
rect 979 17 1013 113
rect 1147 17 1181 113
rect 1315 17 1349 113
rect 1483 17 1517 113
rect 1651 17 1685 113
rect 1819 17 1853 113
rect 1987 17 2021 113
rect 2155 17 2189 113
rect 2323 17 2357 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< labels >>
rlabel locali s 22 215 88 255 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 2392 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 2391 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 2430 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 2392 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1399 51 1433 52 6 X
port 6 nsew signal output
rlabel locali s 1231 51 1265 52 6 X
port 6 nsew signal output
rlabel locali s 1047 51 1097 52 6 X
port 6 nsew signal output
rlabel locali s 2223 52 2289 147 6 X
port 6 nsew signal output
rlabel locali s 2055 52 2121 147 6 X
port 6 nsew signal output
rlabel locali s 1887 52 1953 147 6 X
port 6 nsew signal output
rlabel locali s 1719 52 1785 147 6 X
port 6 nsew signal output
rlabel locali s 1551 52 1617 147 6 X
port 6 nsew signal output
rlabel locali s 1383 52 1449 147 6 X
port 6 nsew signal output
rlabel locali s 1215 52 1281 147 6 X
port 6 nsew signal output
rlabel locali s 1047 52 1113 147 6 X
port 6 nsew signal output
rlabel locali s 1047 147 2375 181 6 X
port 6 nsew signal output
rlabel locali s 2324 181 2375 289 6 X
port 6 nsew signal output
rlabel locali s 1047 289 2375 323 6 X
port 6 nsew signal output
rlabel locali s 2223 323 2289 493 6 X
port 6 nsew signal output
rlabel locali s 2055 323 2121 493 6 X
port 6 nsew signal output
rlabel locali s 1887 323 1953 493 6 X
port 6 nsew signal output
rlabel locali s 1719 323 1785 493 6 X
port 6 nsew signal output
rlabel locali s 1551 323 1617 493 6 X
port 6 nsew signal output
rlabel locali s 1383 323 1449 493 6 X
port 6 nsew signal output
rlabel locali s 1215 323 1281 493 6 X
port 6 nsew signal output
rlabel locali s 1047 323 1113 493 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2392 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3248420
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3230218
<< end >>
