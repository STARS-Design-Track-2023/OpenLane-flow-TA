magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< locali >>
rect 0 1397 746 1431
rect 330 686 364 1151
rect 330 652 459 686
rect 557 652 591 686
rect 212 485 246 551
rect 112 237 146 303
rect 0 -17 746 17
use sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_0  sky130_sram_2kbyte_1rw1r_32x512_8_pdriver_0_0
timestamp 1686671242
transform 1 0 378 0 1 0
box -36 -17 404 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pnand2_0  sky130_sram_2kbyte_1rw1r_32x512_8_pnand2_0_0
timestamp 1686671242
transform 1 0 0 0 1 0
box -36 -17 414 1471
<< labels >>
rlabel locali s 574 669 574 669 4 Z
rlabel locali s 129 270 129 270 4 A
rlabel locali s 229 518 229 518 4 B
rlabel locali s 373 0 373 0 4 gnd
rlabel locali s 373 1414 373 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 746 1414
string GDS_END 396344
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 395202
<< end >>
