magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 1 21 367 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 175 47 205 177
rect 259 47 289 177
<< scpmoshvt >>
rect 79 297 109 497
rect 151 297 181 497
rect 259 357 289 497
<< ndiff >>
rect 27 103 79 177
rect 27 69 35 103
rect 69 69 79 103
rect 27 47 79 69
rect 109 89 175 177
rect 109 55 131 89
rect 165 55 175 89
rect 109 47 175 55
rect 205 112 259 177
rect 205 78 215 112
rect 249 78 259 112
rect 205 47 259 78
rect 289 128 341 177
rect 289 94 299 128
rect 333 94 341 128
rect 289 47 341 94
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 297 151 497
rect 181 485 259 497
rect 181 451 209 485
rect 243 451 259 485
rect 181 417 259 451
rect 181 383 209 417
rect 243 383 259 417
rect 181 357 259 383
rect 289 485 341 497
rect 289 451 299 485
rect 333 451 341 485
rect 289 417 341 451
rect 289 383 299 417
rect 333 383 341 417
rect 289 357 341 383
rect 181 297 231 357
<< ndiffc >>
rect 35 69 69 103
rect 131 55 165 89
rect 215 78 249 112
rect 299 94 333 128
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 209 451 243 485
rect 209 383 243 417
rect 299 451 333 485
rect 299 383 333 417
<< poly >>
rect 79 497 109 523
rect 151 497 181 523
rect 259 497 289 523
rect 259 325 289 357
rect 259 309 347 325
rect 79 265 109 297
rect 38 249 109 265
rect 38 215 48 249
rect 82 215 109 249
rect 38 199 109 215
rect 151 265 181 297
rect 259 275 303 309
rect 337 275 347 309
rect 151 249 207 265
rect 151 215 161 249
rect 195 215 207 249
rect 151 199 207 215
rect 259 259 347 275
rect 79 177 109 199
rect 175 177 205 199
rect 259 177 289 259
rect 79 21 109 47
rect 175 21 205 47
rect 259 21 289 47
<< polycont >>
rect 48 215 82 249
rect 303 275 337 309
rect 161 215 195 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 18 485 82 527
rect 18 451 35 485
rect 69 451 82 485
rect 193 485 259 493
rect 18 417 82 451
rect 18 383 35 417
rect 69 383 82 417
rect 18 349 82 383
rect 18 315 35 349
rect 69 315 82 349
rect 18 299 82 315
rect 118 265 157 475
rect 193 451 209 485
rect 243 451 259 485
rect 193 417 259 451
rect 193 383 209 417
rect 243 383 259 417
rect 193 357 259 383
rect 299 485 350 527
rect 333 451 350 485
rect 299 417 350 451
rect 333 383 350 417
rect 299 367 350 383
rect 193 301 263 357
rect 30 249 82 265
rect 30 215 48 249
rect 30 199 82 215
rect 118 249 195 265
rect 118 215 161 249
rect 118 199 195 215
rect 229 225 263 301
rect 301 309 350 331
rect 301 275 303 309
rect 337 275 350 309
rect 301 259 350 275
rect 229 191 333 225
rect 18 123 261 157
rect 18 103 76 123
rect 18 69 35 103
rect 69 69 76 103
rect 215 112 261 123
rect 18 53 76 69
rect 115 55 131 89
rect 165 55 181 89
rect 249 78 261 112
rect 299 128 333 191
rect 299 78 333 94
rect 215 62 261 78
rect 115 17 181 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 122 425 156 459 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 122 357 156 391 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 122 289 156 323 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 305 289 339 323 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 214 425 248 459 0 FreeSans 400 0 0 0 Y
port 8 nsew signal output
flabel locali s 214 357 248 391 0 FreeSans 400 0 0 0 Y
port 8 nsew signal output
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 o21ai_1
rlabel metal1 s 0 -48 368 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 368 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_END 1275244
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1270526
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 1.840 2.720 
<< end >>
