magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 459 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 182 47 212 177
rect 267 47 297 177
rect 351 47 381 177
<< scpmoshvt >>
rect 79 297 109 497
rect 161 297 191 497
rect 267 297 297 497
rect 351 297 381 497
<< ndiff >>
rect 27 95 79 177
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 127 182 177
rect 109 93 138 127
rect 172 93 182 127
rect 109 47 182 93
rect 212 95 267 177
rect 212 61 223 95
rect 257 61 267 95
rect 212 47 267 61
rect 297 127 351 177
rect 297 93 307 127
rect 341 93 351 127
rect 297 47 351 93
rect 381 95 433 177
rect 381 61 391 95
rect 425 61 433 95
rect 381 47 433 61
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 297 161 497
rect 191 297 267 497
rect 297 297 351 497
rect 381 485 433 497
rect 381 451 391 485
rect 425 451 433 485
rect 381 417 433 451
rect 381 383 391 417
rect 425 383 433 417
rect 381 297 433 383
<< ndiffc >>
rect 35 61 69 95
rect 138 93 172 127
rect 223 61 257 95
rect 307 93 341 127
rect 391 61 425 95
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 391 451 425 485
rect 391 383 425 417
<< poly >>
rect 79 497 109 523
rect 161 497 191 523
rect 267 497 297 523
rect 351 497 381 523
rect 79 265 109 297
rect 161 265 191 297
rect 267 265 297 297
rect 351 265 381 297
rect 21 249 109 265
rect 21 215 33 249
rect 67 215 109 249
rect 21 199 109 215
rect 159 249 213 265
rect 159 215 169 249
rect 203 215 213 249
rect 159 199 213 215
rect 255 249 309 265
rect 255 215 265 249
rect 299 215 309 249
rect 255 199 309 215
rect 351 249 439 265
rect 351 215 395 249
rect 429 215 439 249
rect 351 199 439 215
rect 79 177 109 199
rect 182 177 212 199
rect 267 177 297 199
rect 351 177 381 199
rect 79 21 109 47
rect 182 21 212 47
rect 267 21 297 47
rect 351 21 381 47
<< polycont >>
rect 33 215 67 249
rect 169 215 203 249
rect 265 215 299 249
rect 395 215 429 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 18 485 85 490
rect 18 451 35 485
rect 69 451 85 485
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 18 349 85 383
rect 18 315 35 349
rect 69 333 85 349
rect 69 315 135 333
rect 206 323 257 490
rect 18 299 135 315
rect 17 249 67 265
rect 17 215 33 249
rect 17 149 67 215
rect 101 165 135 299
rect 169 283 257 323
rect 169 249 215 283
rect 291 249 339 490
rect 391 485 443 527
rect 425 451 443 485
rect 391 417 443 451
rect 425 383 443 417
rect 391 367 443 383
rect 203 215 215 249
rect 249 215 265 249
rect 299 215 339 249
rect 391 249 443 333
rect 391 215 395 249
rect 429 215 443 249
rect 169 199 215 215
rect 101 131 341 165
rect 391 131 443 215
rect 101 129 172 131
rect 119 127 172 129
rect 17 95 69 115
rect 17 61 35 95
rect 119 93 138 127
rect 307 127 341 131
rect 119 77 172 93
rect 207 95 273 97
rect 17 17 69 61
rect 207 61 223 95
rect 257 61 273 95
rect 307 77 341 93
rect 375 95 441 97
rect 207 17 273 61
rect 375 61 391 95
rect 425 61 441 95
rect 375 17 441 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 29 153 63 187 0 FreeSans 400 0 0 0 D
port 4 nsew signal input
flabel locali s 213 289 247 323 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 28 221 62 255 0 FreeSans 400 0 0 0 D
port 4 nsew signal input
flabel locali s 30 425 64 459 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 397 153 431 187 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 305 357 339 391 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor4_1
rlabel metal1 s 0 -48 460 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 1132892
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1128172
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 2.300 0.000 
<< end >>
