magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1451 203
rect 29 -17 63 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 419 47 449 177
rect 503 47 533 177
rect 587 47 617 177
rect 671 47 701 177
rect 755 47 785 177
rect 839 47 869 177
rect 923 47 953 177
rect 1007 47 1037 177
rect 1091 47 1121 177
rect 1175 47 1205 177
rect 1259 47 1289 177
rect 1343 47 1373 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 419 297 449 497
rect 503 297 533 497
rect 587 297 617 497
rect 671 297 701 497
rect 755 297 785 497
rect 839 297 869 497
rect 923 297 953 497
rect 1007 297 1037 497
rect 1091 297 1121 497
rect 1175 297 1205 497
rect 1259 297 1289 497
rect 1343 297 1373 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 95 335 129
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 95 419 177
rect 365 61 375 95
rect 409 61 419 95
rect 365 47 419 61
rect 449 163 503 177
rect 449 129 459 163
rect 493 129 503 163
rect 449 95 503 129
rect 449 61 459 95
rect 493 61 503 95
rect 449 47 503 61
rect 533 95 587 177
rect 533 61 543 95
rect 577 61 587 95
rect 533 47 587 61
rect 617 163 671 177
rect 617 129 627 163
rect 661 129 671 163
rect 617 95 671 129
rect 617 61 627 95
rect 661 61 671 95
rect 617 47 671 61
rect 701 95 755 177
rect 701 61 711 95
rect 745 61 755 95
rect 701 47 755 61
rect 785 163 839 177
rect 785 129 795 163
rect 829 129 839 163
rect 785 95 839 129
rect 785 61 795 95
rect 829 61 839 95
rect 785 47 839 61
rect 869 95 923 177
rect 869 61 879 95
rect 913 61 923 95
rect 869 47 923 61
rect 953 163 1007 177
rect 953 129 963 163
rect 997 129 1007 163
rect 953 95 1007 129
rect 953 61 963 95
rect 997 61 1007 95
rect 953 47 1007 61
rect 1037 95 1091 177
rect 1037 61 1047 95
rect 1081 61 1091 95
rect 1037 47 1091 61
rect 1121 163 1175 177
rect 1121 129 1131 163
rect 1165 129 1175 163
rect 1121 95 1175 129
rect 1121 61 1131 95
rect 1165 61 1175 95
rect 1121 47 1175 61
rect 1205 95 1259 177
rect 1205 61 1215 95
rect 1249 61 1259 95
rect 1205 47 1259 61
rect 1289 163 1343 177
rect 1289 129 1299 163
rect 1333 129 1343 163
rect 1289 95 1343 129
rect 1289 61 1299 95
rect 1333 61 1343 95
rect 1289 47 1343 61
rect 1373 95 1425 177
rect 1373 61 1383 95
rect 1417 61 1425 95
rect 1373 47 1425 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 485 167 497
rect 113 451 123 485
rect 157 451 167 485
rect 113 417 167 451
rect 113 383 123 417
rect 157 383 167 417
rect 113 297 167 383
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 341 251 375
rect 197 307 207 341
rect 241 307 251 341
rect 197 297 251 307
rect 281 485 335 497
rect 281 451 291 485
rect 325 451 335 485
rect 281 417 335 451
rect 281 383 291 417
rect 325 383 335 417
rect 281 297 335 383
rect 365 477 419 497
rect 365 443 375 477
rect 409 443 419 477
rect 365 409 419 443
rect 365 375 375 409
rect 409 375 419 409
rect 365 341 419 375
rect 365 307 375 341
rect 409 307 419 341
rect 365 297 419 307
rect 449 485 503 497
rect 449 451 459 485
rect 493 451 503 485
rect 449 417 503 451
rect 449 383 459 417
rect 493 383 503 417
rect 449 297 503 383
rect 533 477 587 497
rect 533 443 543 477
rect 577 443 587 477
rect 533 409 587 443
rect 533 375 543 409
rect 577 375 587 409
rect 533 341 587 375
rect 533 307 543 341
rect 577 307 587 341
rect 533 297 587 307
rect 617 485 671 497
rect 617 451 627 485
rect 661 451 671 485
rect 617 417 671 451
rect 617 383 627 417
rect 661 383 671 417
rect 617 297 671 383
rect 701 477 755 497
rect 701 443 711 477
rect 745 443 755 477
rect 701 409 755 443
rect 701 375 711 409
rect 745 375 755 409
rect 701 341 755 375
rect 701 307 711 341
rect 745 307 755 341
rect 701 297 755 307
rect 785 409 839 497
rect 785 375 795 409
rect 829 375 839 409
rect 785 341 839 375
rect 785 307 795 341
rect 829 307 839 341
rect 785 297 839 307
rect 869 477 923 497
rect 869 443 879 477
rect 913 443 923 477
rect 869 409 923 443
rect 869 375 879 409
rect 913 375 923 409
rect 869 297 923 375
rect 953 409 1007 497
rect 953 375 963 409
rect 997 375 1007 409
rect 953 341 1007 375
rect 953 307 963 341
rect 997 307 1007 341
rect 953 297 1007 307
rect 1037 477 1091 497
rect 1037 443 1047 477
rect 1081 443 1091 477
rect 1037 409 1091 443
rect 1037 375 1047 409
rect 1081 375 1091 409
rect 1037 297 1091 375
rect 1121 409 1175 497
rect 1121 375 1131 409
rect 1165 375 1175 409
rect 1121 341 1175 375
rect 1121 307 1131 341
rect 1165 307 1175 341
rect 1121 297 1175 307
rect 1205 477 1259 497
rect 1205 443 1215 477
rect 1249 443 1259 477
rect 1205 409 1259 443
rect 1205 375 1215 409
rect 1249 375 1259 409
rect 1205 297 1259 375
rect 1289 409 1343 497
rect 1289 375 1299 409
rect 1333 375 1343 409
rect 1289 341 1343 375
rect 1289 307 1299 341
rect 1333 307 1343 341
rect 1289 297 1343 307
rect 1373 477 1427 497
rect 1373 443 1383 477
rect 1417 443 1427 477
rect 1373 409 1427 443
rect 1373 375 1383 409
rect 1417 375 1427 409
rect 1373 297 1427 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 61 241 95
rect 291 129 325 163
rect 291 61 325 95
rect 375 61 409 95
rect 459 129 493 163
rect 459 61 493 95
rect 543 61 577 95
rect 627 129 661 163
rect 627 61 661 95
rect 711 61 745 95
rect 795 129 829 163
rect 795 61 829 95
rect 879 61 913 95
rect 963 129 997 163
rect 963 61 997 95
rect 1047 61 1081 95
rect 1131 129 1165 163
rect 1131 61 1165 95
rect 1215 61 1249 95
rect 1299 129 1333 163
rect 1299 61 1333 95
rect 1383 61 1417 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 451 157 485
rect 123 383 157 417
rect 207 443 241 477
rect 207 375 241 409
rect 207 307 241 341
rect 291 451 325 485
rect 291 383 325 417
rect 375 443 409 477
rect 375 375 409 409
rect 375 307 409 341
rect 459 451 493 485
rect 459 383 493 417
rect 543 443 577 477
rect 543 375 577 409
rect 543 307 577 341
rect 627 451 661 485
rect 627 383 661 417
rect 711 443 745 477
rect 711 375 745 409
rect 711 307 745 341
rect 795 375 829 409
rect 795 307 829 341
rect 879 443 913 477
rect 879 375 913 409
rect 963 375 997 409
rect 963 307 997 341
rect 1047 443 1081 477
rect 1047 375 1081 409
rect 1131 375 1165 409
rect 1131 307 1165 341
rect 1215 443 1249 477
rect 1215 375 1249 409
rect 1299 375 1333 409
rect 1299 307 1333 341
rect 1383 443 1417 477
rect 1383 375 1417 409
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 419 497 449 523
rect 503 497 533 523
rect 587 497 617 523
rect 671 497 701 523
rect 755 497 785 523
rect 839 497 869 523
rect 923 497 953 523
rect 1007 497 1037 523
rect 1091 497 1121 523
rect 1175 497 1205 523
rect 1259 497 1289 523
rect 1343 497 1373 523
rect 83 265 113 297
rect 167 265 197 297
rect 251 265 281 297
rect 335 265 365 297
rect 419 265 449 297
rect 503 265 533 297
rect 587 265 617 297
rect 671 265 701 297
rect 83 249 701 265
rect 83 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 375 249
rect 409 215 443 249
rect 477 215 511 249
rect 545 215 579 249
rect 613 215 647 249
rect 681 215 701 249
rect 83 199 701 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 177 281 199
rect 335 177 365 199
rect 419 177 449 199
rect 503 177 533 199
rect 587 177 617 199
rect 671 177 701 199
rect 755 265 785 297
rect 839 265 869 297
rect 923 265 953 297
rect 1007 265 1037 297
rect 1091 265 1121 297
rect 1175 265 1205 297
rect 1259 265 1289 297
rect 1343 265 1373 297
rect 755 249 1373 265
rect 755 215 778 249
rect 812 215 846 249
rect 880 215 914 249
rect 948 215 982 249
rect 1016 215 1050 249
rect 1084 215 1118 249
rect 1152 215 1186 249
rect 1220 215 1254 249
rect 1288 215 1373 249
rect 755 199 1373 215
rect 755 177 785 199
rect 839 177 869 199
rect 923 177 953 199
rect 1007 177 1037 199
rect 1091 177 1121 199
rect 1175 177 1205 199
rect 1259 177 1289 199
rect 1343 177 1373 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 419 21 449 47
rect 503 21 533 47
rect 587 21 617 47
rect 671 21 701 47
rect 755 21 785 47
rect 839 21 869 47
rect 923 21 953 47
rect 1007 21 1037 47
rect 1091 21 1121 47
rect 1175 21 1205 47
rect 1259 21 1289 47
rect 1343 21 1373 47
<< polycont >>
rect 103 215 137 249
rect 171 215 205 249
rect 239 215 273 249
rect 307 215 341 249
rect 375 215 409 249
rect 443 215 477 249
rect 511 215 545 249
rect 579 215 613 249
rect 647 215 681 249
rect 778 215 812 249
rect 846 215 880 249
rect 914 215 948 249
rect 982 215 1016 249
rect 1050 215 1084 249
rect 1118 215 1152 249
rect 1186 215 1220 249
rect 1254 215 1288 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 18 477 81 493
rect 18 443 39 477
rect 73 443 81 477
rect 18 409 81 443
rect 18 375 39 409
rect 73 375 81 409
rect 18 341 81 375
rect 115 485 165 527
rect 115 451 123 485
rect 157 451 165 485
rect 115 417 165 451
rect 115 383 123 417
rect 157 383 165 417
rect 115 367 165 383
rect 199 477 249 493
rect 199 443 207 477
rect 241 443 249 477
rect 199 409 249 443
rect 199 375 207 409
rect 241 375 249 409
rect 18 307 39 341
rect 73 333 81 341
rect 199 341 249 375
rect 283 485 333 527
rect 283 451 291 485
rect 325 451 333 485
rect 283 417 333 451
rect 283 383 291 417
rect 325 383 333 417
rect 283 367 333 383
rect 367 477 417 493
rect 367 443 375 477
rect 409 443 417 477
rect 367 409 417 443
rect 367 375 375 409
rect 409 375 417 409
rect 199 333 207 341
rect 73 307 207 333
rect 241 333 249 341
rect 367 341 417 375
rect 451 485 501 527
rect 451 451 459 485
rect 493 451 501 485
rect 451 417 501 451
rect 451 383 459 417
rect 493 383 501 417
rect 451 367 501 383
rect 535 477 585 493
rect 535 443 543 477
rect 577 443 585 477
rect 535 409 585 443
rect 535 375 543 409
rect 577 375 585 409
rect 367 333 375 341
rect 241 307 375 333
rect 409 333 417 341
rect 535 341 585 375
rect 619 485 669 527
rect 619 451 627 485
rect 661 451 669 485
rect 619 417 669 451
rect 619 383 627 417
rect 661 383 669 417
rect 619 367 669 383
rect 703 477 1425 493
rect 703 443 711 477
rect 745 459 879 477
rect 745 443 753 459
rect 703 409 753 443
rect 871 443 879 459
rect 913 459 1047 477
rect 913 443 921 459
rect 703 375 711 409
rect 745 375 753 409
rect 535 333 543 341
rect 409 307 543 333
rect 577 333 585 341
rect 703 341 753 375
rect 703 333 711 341
rect 577 307 711 333
rect 745 307 753 341
rect 18 291 753 307
rect 787 409 837 425
rect 787 375 795 409
rect 829 375 837 409
rect 787 341 837 375
rect 871 409 921 443
rect 1039 443 1047 459
rect 1081 459 1215 477
rect 1081 443 1089 459
rect 871 375 879 409
rect 913 375 921 409
rect 871 357 921 375
rect 955 409 1005 425
rect 955 375 963 409
rect 997 375 1005 409
rect 787 307 795 341
rect 829 323 837 341
rect 955 341 1005 375
rect 1039 409 1089 443
rect 1207 443 1215 459
rect 1249 459 1383 477
rect 1249 443 1257 459
rect 1039 375 1047 409
rect 1081 375 1089 409
rect 1039 357 1089 375
rect 1123 409 1173 425
rect 1123 375 1131 409
rect 1165 375 1173 409
rect 955 323 963 341
rect 829 307 963 323
rect 997 323 1005 341
rect 1123 341 1173 375
rect 1207 409 1257 443
rect 1375 443 1383 459
rect 1417 443 1425 477
rect 1207 375 1215 409
rect 1249 375 1257 409
rect 1207 357 1257 375
rect 1291 409 1341 425
rect 1291 375 1299 409
rect 1333 375 1341 409
rect 1123 323 1131 341
rect 997 307 1131 323
rect 1165 323 1173 341
rect 1291 341 1341 375
rect 1375 409 1425 443
rect 1375 375 1383 409
rect 1417 375 1425 409
rect 1375 357 1425 375
rect 1291 323 1299 341
rect 1165 307 1299 323
rect 1333 323 1341 341
rect 1333 307 1455 323
rect 787 289 1455 307
rect 72 249 706 255
rect 72 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 375 249
rect 409 215 443 249
rect 477 215 511 249
rect 545 215 579 249
rect 613 215 647 249
rect 681 215 706 249
rect 760 249 1308 255
rect 760 215 778 249
rect 812 215 846 249
rect 880 215 914 249
rect 948 215 982 249
rect 1016 215 1050 249
rect 1084 215 1118 249
rect 1152 215 1186 249
rect 1220 215 1254 249
rect 1288 215 1308 249
rect 1342 181 1455 289
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 1455 181
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 107 95 173 129
rect 275 129 291 145
rect 325 145 459 163
rect 325 129 341 145
rect 107 61 123 95
rect 157 61 173 95
rect 107 51 173 61
rect 207 95 241 111
rect 207 17 241 61
rect 275 95 341 129
rect 443 129 459 145
rect 493 145 627 163
rect 493 129 509 145
rect 275 61 291 95
rect 325 61 341 95
rect 275 51 341 61
rect 375 95 409 111
rect 375 17 409 61
rect 443 95 509 129
rect 611 129 627 145
rect 661 145 795 163
rect 661 129 677 145
rect 443 61 459 95
rect 493 61 509 95
rect 443 51 509 61
rect 543 95 577 111
rect 543 17 577 61
rect 611 95 677 129
rect 779 129 795 145
rect 829 145 963 163
rect 829 129 845 145
rect 611 61 627 95
rect 661 61 677 95
rect 611 51 677 61
rect 711 95 745 111
rect 711 17 745 61
rect 779 95 845 129
rect 947 129 963 145
rect 997 145 1131 163
rect 997 129 1013 145
rect 779 61 795 95
rect 829 61 845 95
rect 779 51 845 61
rect 879 95 913 111
rect 879 17 913 61
rect 947 95 1013 129
rect 1115 129 1131 145
rect 1165 145 1299 163
rect 1165 129 1181 145
rect 947 61 963 95
rect 997 61 1013 95
rect 947 51 1013 61
rect 1047 95 1081 111
rect 1047 17 1081 61
rect 1115 95 1181 129
rect 1283 129 1299 145
rect 1333 145 1455 163
rect 1333 129 1349 145
rect 1115 61 1131 95
rect 1165 61 1181 95
rect 1115 51 1181 61
rect 1215 95 1249 111
rect 1215 17 1249 61
rect 1283 95 1349 129
rect 1283 61 1299 95
rect 1333 61 1349 95
rect 1283 51 1349 61
rect 1383 95 1441 111
rect 1417 61 1441 95
rect 1383 17 1441 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel locali s 1409 289 1443 323 0 FreeSans 400 0 0 0 Y
port 7 nsew signal output
flabel locali s 121 221 155 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor2_8
rlabel metal1 s 0 -48 1472 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1472 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_END 1980998
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1969600
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 36.800 0.000 
<< end >>
