magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__dfl1sd__example_5595914180872  sky130_fd_pr__dfl1sd__example_5595914180872_0
timestamp 1686671242
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180872  sky130_fd_pr__dfl1sd__example_5595914180872_1
timestamp 1686671242
transform 1 0 120 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 40245314
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 40244264
<< end >>
