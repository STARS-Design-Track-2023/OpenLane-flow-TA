magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_0
timestamp 1686671242
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_1
timestamp 1686671242
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_2
timestamp 1686671242
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_3
timestamp 1686671242
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_4
timestamp 1686671242
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_5
timestamp 1686671242
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_6
timestamp 1686671242
transform 1 0 880 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_7
timestamp 1686671242
transform 1 0 1036 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_8
timestamp 1686671242
transform 1 0 1192 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_9
timestamp 1686671242
transform 1 0 1348 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_10
timestamp 1686671242
transform 1 0 1504 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_11
timestamp 1686671242
transform 1 0 1660 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_12
timestamp 1686671242
transform 1 0 1816 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_13
timestamp 1686671242
transform 1 0 1972 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_14
timestamp 1686671242
transform 1 0 2128 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 8080164
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8072500
<< end >>
