magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 63 21 1745 203
rect 29 -17 63 17
<< scnmos >>
rect 141 47 171 177
rect 225 47 255 177
rect 377 47 407 177
rect 461 47 491 177
rect 545 47 575 177
rect 629 47 659 177
rect 713 47 743 177
rect 797 47 827 177
rect 881 47 911 177
rect 965 47 995 177
rect 1049 47 1079 177
rect 1133 47 1163 177
rect 1217 47 1247 177
rect 1301 47 1331 177
rect 1385 47 1415 177
rect 1469 47 1499 177
rect 1553 47 1583 177
rect 1637 47 1667 177
<< scpmoshvt >>
rect 93 297 123 497
rect 177 297 207 497
rect 377 297 407 497
rect 461 297 491 497
rect 545 297 575 497
rect 629 297 659 497
rect 713 297 743 497
rect 797 297 827 497
rect 881 297 911 497
rect 965 297 995 497
rect 1049 297 1079 497
rect 1133 297 1163 497
rect 1217 297 1247 497
rect 1301 297 1331 497
rect 1385 297 1415 497
rect 1469 297 1499 497
rect 1553 297 1583 497
rect 1637 297 1667 497
<< ndiff >>
rect 89 163 141 177
rect 89 129 97 163
rect 131 129 141 163
rect 89 95 141 129
rect 89 61 97 95
rect 131 61 141 95
rect 89 47 141 61
rect 171 163 225 177
rect 171 129 181 163
rect 215 129 225 163
rect 171 95 225 129
rect 171 61 181 95
rect 215 61 225 95
rect 171 47 225 61
rect 255 163 377 177
rect 255 61 265 163
rect 367 61 377 163
rect 255 47 377 61
rect 407 163 461 177
rect 407 129 417 163
rect 451 129 461 163
rect 407 95 461 129
rect 407 61 417 95
rect 451 61 461 95
rect 407 47 461 61
rect 491 95 545 177
rect 491 61 501 95
rect 535 61 545 95
rect 491 47 545 61
rect 575 163 629 177
rect 575 129 585 163
rect 619 129 629 163
rect 575 95 629 129
rect 575 61 585 95
rect 619 61 629 95
rect 575 47 629 61
rect 659 95 713 177
rect 659 61 669 95
rect 703 61 713 95
rect 659 47 713 61
rect 743 163 797 177
rect 743 129 753 163
rect 787 129 797 163
rect 743 95 797 129
rect 743 61 753 95
rect 787 61 797 95
rect 743 47 797 61
rect 827 95 881 177
rect 827 61 837 95
rect 871 61 881 95
rect 827 47 881 61
rect 911 163 965 177
rect 911 129 921 163
rect 955 129 965 163
rect 911 95 965 129
rect 911 61 921 95
rect 955 61 965 95
rect 911 47 965 61
rect 995 95 1049 177
rect 995 61 1005 95
rect 1039 61 1049 95
rect 995 47 1049 61
rect 1079 163 1133 177
rect 1079 129 1089 163
rect 1123 129 1133 163
rect 1079 95 1133 129
rect 1079 61 1089 95
rect 1123 61 1133 95
rect 1079 47 1133 61
rect 1163 95 1217 177
rect 1163 61 1173 95
rect 1207 61 1217 95
rect 1163 47 1217 61
rect 1247 163 1301 177
rect 1247 129 1257 163
rect 1291 129 1301 163
rect 1247 95 1301 129
rect 1247 61 1257 95
rect 1291 61 1301 95
rect 1247 47 1301 61
rect 1331 95 1385 177
rect 1331 61 1341 95
rect 1375 61 1385 95
rect 1331 47 1385 61
rect 1415 163 1469 177
rect 1415 129 1425 163
rect 1459 129 1469 163
rect 1415 95 1469 129
rect 1415 61 1425 95
rect 1459 61 1469 95
rect 1415 47 1469 61
rect 1499 95 1553 177
rect 1499 61 1509 95
rect 1543 61 1553 95
rect 1499 47 1553 61
rect 1583 163 1637 177
rect 1583 129 1593 163
rect 1627 129 1637 163
rect 1583 95 1637 129
rect 1583 61 1593 95
rect 1627 61 1637 95
rect 1583 47 1637 61
rect 1667 95 1719 177
rect 1667 61 1677 95
rect 1711 61 1719 95
rect 1667 47 1719 61
<< pdiff >>
rect 41 485 93 497
rect 41 451 49 485
rect 83 451 93 485
rect 41 415 93 451
rect 41 381 49 415
rect 83 381 93 415
rect 41 345 93 381
rect 41 311 49 345
rect 83 311 93 345
rect 41 297 93 311
rect 123 477 177 497
rect 123 443 133 477
rect 167 443 177 477
rect 123 409 177 443
rect 123 375 133 409
rect 167 375 177 409
rect 123 341 177 375
rect 123 307 133 341
rect 167 307 177 341
rect 123 297 177 307
rect 207 485 263 497
rect 207 451 217 485
rect 251 451 263 485
rect 207 415 263 451
rect 207 381 217 415
rect 251 381 263 415
rect 207 345 263 381
rect 207 311 217 345
rect 251 311 263 345
rect 207 297 263 311
rect 321 477 377 497
rect 321 443 333 477
rect 367 443 377 477
rect 321 409 377 443
rect 321 375 333 409
rect 367 375 377 409
rect 321 341 377 375
rect 321 307 333 341
rect 367 307 377 341
rect 321 297 377 307
rect 407 485 461 497
rect 407 451 417 485
rect 451 451 461 485
rect 407 417 461 451
rect 407 383 417 417
rect 451 383 461 417
rect 407 297 461 383
rect 491 477 545 497
rect 491 443 501 477
rect 535 443 545 477
rect 491 409 545 443
rect 491 375 501 409
rect 535 375 545 409
rect 491 341 545 375
rect 491 307 501 341
rect 535 307 545 341
rect 491 297 545 307
rect 575 485 629 497
rect 575 451 585 485
rect 619 451 629 485
rect 575 417 629 451
rect 575 383 585 417
rect 619 383 629 417
rect 575 297 629 383
rect 659 477 713 497
rect 659 443 669 477
rect 703 443 713 477
rect 659 409 713 443
rect 659 375 669 409
rect 703 375 713 409
rect 659 341 713 375
rect 659 307 669 341
rect 703 307 713 341
rect 659 297 713 307
rect 743 485 797 497
rect 743 451 753 485
rect 787 451 797 485
rect 743 417 797 451
rect 743 383 753 417
rect 787 383 797 417
rect 743 297 797 383
rect 827 477 881 497
rect 827 443 837 477
rect 871 443 881 477
rect 827 409 881 443
rect 827 375 837 409
rect 871 375 881 409
rect 827 341 881 375
rect 827 307 837 341
rect 871 307 881 341
rect 827 297 881 307
rect 911 485 965 497
rect 911 451 921 485
rect 955 451 965 485
rect 911 417 965 451
rect 911 383 921 417
rect 955 383 965 417
rect 911 297 965 383
rect 995 477 1049 497
rect 995 443 1005 477
rect 1039 443 1049 477
rect 995 409 1049 443
rect 995 375 1005 409
rect 1039 375 1049 409
rect 995 341 1049 375
rect 995 307 1005 341
rect 1039 307 1049 341
rect 995 297 1049 307
rect 1079 409 1133 497
rect 1079 375 1089 409
rect 1123 375 1133 409
rect 1079 341 1133 375
rect 1079 307 1089 341
rect 1123 307 1133 341
rect 1079 297 1133 307
rect 1163 477 1217 497
rect 1163 443 1173 477
rect 1207 443 1217 477
rect 1163 409 1217 443
rect 1163 375 1173 409
rect 1207 375 1217 409
rect 1163 297 1217 375
rect 1247 409 1301 497
rect 1247 375 1257 409
rect 1291 375 1301 409
rect 1247 341 1301 375
rect 1247 307 1257 341
rect 1291 307 1301 341
rect 1247 297 1301 307
rect 1331 477 1385 497
rect 1331 443 1341 477
rect 1375 443 1385 477
rect 1331 409 1385 443
rect 1331 375 1341 409
rect 1375 375 1385 409
rect 1331 297 1385 375
rect 1415 409 1469 497
rect 1415 375 1425 409
rect 1459 375 1469 409
rect 1415 341 1469 375
rect 1415 307 1425 341
rect 1459 307 1469 341
rect 1415 297 1469 307
rect 1499 477 1553 497
rect 1499 443 1509 477
rect 1543 443 1553 477
rect 1499 409 1553 443
rect 1499 375 1509 409
rect 1543 375 1553 409
rect 1499 297 1553 375
rect 1583 409 1637 497
rect 1583 375 1593 409
rect 1627 375 1637 409
rect 1583 341 1637 375
rect 1583 307 1593 341
rect 1627 307 1637 341
rect 1583 297 1637 307
rect 1667 477 1721 497
rect 1667 443 1677 477
rect 1711 443 1721 477
rect 1667 409 1721 443
rect 1667 375 1677 409
rect 1711 375 1721 409
rect 1667 297 1721 375
<< ndiffc >>
rect 97 129 131 163
rect 97 61 131 95
rect 181 129 215 163
rect 181 61 215 95
rect 265 61 367 163
rect 417 129 451 163
rect 417 61 451 95
rect 501 61 535 95
rect 585 129 619 163
rect 585 61 619 95
rect 669 61 703 95
rect 753 129 787 163
rect 753 61 787 95
rect 837 61 871 95
rect 921 129 955 163
rect 921 61 955 95
rect 1005 61 1039 95
rect 1089 129 1123 163
rect 1089 61 1123 95
rect 1173 61 1207 95
rect 1257 129 1291 163
rect 1257 61 1291 95
rect 1341 61 1375 95
rect 1425 129 1459 163
rect 1425 61 1459 95
rect 1509 61 1543 95
rect 1593 129 1627 163
rect 1593 61 1627 95
rect 1677 61 1711 95
<< pdiffc >>
rect 49 451 83 485
rect 49 381 83 415
rect 49 311 83 345
rect 133 443 167 477
rect 133 375 167 409
rect 133 307 167 341
rect 217 451 251 485
rect 217 381 251 415
rect 217 311 251 345
rect 333 443 367 477
rect 333 375 367 409
rect 333 307 367 341
rect 417 451 451 485
rect 417 383 451 417
rect 501 443 535 477
rect 501 375 535 409
rect 501 307 535 341
rect 585 451 619 485
rect 585 383 619 417
rect 669 443 703 477
rect 669 375 703 409
rect 669 307 703 341
rect 753 451 787 485
rect 753 383 787 417
rect 837 443 871 477
rect 837 375 871 409
rect 837 307 871 341
rect 921 451 955 485
rect 921 383 955 417
rect 1005 443 1039 477
rect 1005 375 1039 409
rect 1005 307 1039 341
rect 1089 375 1123 409
rect 1089 307 1123 341
rect 1173 443 1207 477
rect 1173 375 1207 409
rect 1257 375 1291 409
rect 1257 307 1291 341
rect 1341 443 1375 477
rect 1341 375 1375 409
rect 1425 375 1459 409
rect 1425 307 1459 341
rect 1509 443 1543 477
rect 1509 375 1543 409
rect 1593 375 1627 409
rect 1593 307 1627 341
rect 1677 443 1711 477
rect 1677 375 1711 409
<< poly >>
rect 93 497 123 523
rect 177 497 207 523
rect 377 497 407 523
rect 461 497 491 523
rect 545 497 575 523
rect 629 497 659 523
rect 713 497 743 523
rect 797 497 827 523
rect 881 497 911 523
rect 965 497 995 523
rect 1049 497 1079 523
rect 1133 497 1163 523
rect 1217 497 1247 523
rect 1301 497 1331 523
rect 1385 497 1415 523
rect 1469 497 1499 523
rect 1553 497 1583 523
rect 1637 497 1667 523
rect 93 265 123 297
rect 177 265 207 297
rect 377 265 407 297
rect 461 265 491 297
rect 545 265 575 297
rect 629 265 659 297
rect 713 265 743 297
rect 797 265 827 297
rect 881 265 911 297
rect 965 265 995 297
rect 35 249 255 265
rect 35 215 55 249
rect 89 215 255 249
rect 35 199 255 215
rect 141 177 171 199
rect 225 177 255 199
rect 377 249 995 265
rect 377 215 397 249
rect 431 215 465 249
rect 499 215 533 249
rect 567 215 601 249
rect 635 215 669 249
rect 703 215 737 249
rect 771 215 805 249
rect 839 215 873 249
rect 907 215 941 249
rect 975 215 995 249
rect 377 199 995 215
rect 377 177 407 199
rect 461 177 491 199
rect 545 177 575 199
rect 629 177 659 199
rect 713 177 743 199
rect 797 177 827 199
rect 881 177 911 199
rect 965 177 995 199
rect 1049 265 1079 297
rect 1133 265 1163 297
rect 1217 265 1247 297
rect 1301 265 1331 297
rect 1385 265 1415 297
rect 1469 265 1499 297
rect 1553 265 1583 297
rect 1637 265 1667 297
rect 1049 249 1667 265
rect 1049 215 1072 249
rect 1106 215 1140 249
rect 1174 215 1208 249
rect 1242 215 1276 249
rect 1310 215 1344 249
rect 1378 215 1412 249
rect 1446 215 1480 249
rect 1514 215 1548 249
rect 1582 215 1667 249
rect 1049 199 1667 215
rect 1049 177 1079 199
rect 1133 177 1163 199
rect 1217 177 1247 199
rect 1301 177 1331 199
rect 1385 177 1415 199
rect 1469 177 1499 199
rect 1553 177 1583 199
rect 1637 177 1667 199
rect 141 21 171 47
rect 225 21 255 47
rect 377 21 407 47
rect 461 21 491 47
rect 545 21 575 47
rect 629 21 659 47
rect 713 21 743 47
rect 797 21 827 47
rect 881 21 911 47
rect 965 21 995 47
rect 1049 21 1079 47
rect 1133 21 1163 47
rect 1217 21 1247 47
rect 1301 21 1331 47
rect 1385 21 1415 47
rect 1469 21 1499 47
rect 1553 21 1583 47
rect 1637 21 1667 47
<< polycont >>
rect 55 215 89 249
rect 397 215 431 249
rect 465 215 499 249
rect 533 215 567 249
rect 601 215 635 249
rect 669 215 703 249
rect 737 215 771 249
rect 805 215 839 249
rect 873 215 907 249
rect 941 215 975 249
rect 1072 215 1106 249
rect 1140 215 1174 249
rect 1208 215 1242 249
rect 1276 215 1310 249
rect 1344 215 1378 249
rect 1412 215 1446 249
rect 1480 215 1514 249
rect 1548 215 1582 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 39 485 83 527
rect 39 451 49 485
rect 39 415 83 451
rect 39 381 49 415
rect 39 345 83 381
rect 39 311 49 345
rect 39 291 83 311
rect 117 477 183 493
rect 117 443 133 477
rect 167 443 183 477
rect 117 409 183 443
rect 117 375 133 409
rect 167 375 183 409
rect 117 341 183 375
rect 117 307 133 341
rect 167 307 183 341
rect 117 291 183 307
rect 217 485 266 527
rect 251 451 266 485
rect 217 415 266 451
rect 251 381 266 415
rect 217 345 266 381
rect 251 311 266 345
rect 217 291 266 311
rect 311 477 375 493
rect 311 443 333 477
rect 367 443 375 477
rect 311 409 375 443
rect 311 375 333 409
rect 367 375 375 409
rect 311 341 375 375
rect 409 485 459 527
rect 409 451 417 485
rect 451 451 459 485
rect 409 417 459 451
rect 409 383 417 417
rect 451 383 459 417
rect 409 367 459 383
rect 493 477 543 493
rect 493 443 501 477
rect 535 443 543 477
rect 493 409 543 443
rect 493 375 501 409
rect 535 375 543 409
rect 311 307 333 341
rect 367 333 375 341
rect 493 341 543 375
rect 577 485 627 527
rect 577 451 585 485
rect 619 451 627 485
rect 577 417 627 451
rect 577 383 585 417
rect 619 383 627 417
rect 577 367 627 383
rect 661 477 711 493
rect 661 443 669 477
rect 703 443 711 477
rect 661 409 711 443
rect 661 375 669 409
rect 703 375 711 409
rect 493 333 501 341
rect 367 307 501 333
rect 535 333 543 341
rect 661 341 711 375
rect 745 485 795 527
rect 745 451 753 485
rect 787 451 795 485
rect 745 417 795 451
rect 745 383 753 417
rect 787 383 795 417
rect 745 367 795 383
rect 829 477 879 493
rect 829 443 837 477
rect 871 443 879 477
rect 829 409 879 443
rect 829 375 837 409
rect 871 375 879 409
rect 661 333 669 341
rect 535 307 669 333
rect 703 333 711 341
rect 829 341 879 375
rect 913 485 963 527
rect 913 451 921 485
rect 955 451 963 485
rect 913 417 963 451
rect 913 383 921 417
rect 955 383 963 417
rect 913 367 963 383
rect 997 477 1719 493
rect 997 443 1005 477
rect 1039 459 1173 477
rect 1039 443 1047 459
rect 997 409 1047 443
rect 1165 443 1173 459
rect 1207 459 1341 477
rect 1207 443 1215 459
rect 997 375 1005 409
rect 1039 375 1047 409
rect 829 333 837 341
rect 703 307 837 333
rect 871 333 879 341
rect 997 341 1047 375
rect 997 333 1005 341
rect 871 307 1005 333
rect 1039 307 1047 341
rect 311 291 1047 307
rect 1081 409 1131 425
rect 1081 375 1089 409
rect 1123 375 1131 409
rect 1081 341 1131 375
rect 1165 409 1215 443
rect 1333 443 1341 459
rect 1375 459 1509 477
rect 1375 443 1383 459
rect 1165 375 1173 409
rect 1207 375 1215 409
rect 1165 357 1215 375
rect 1249 409 1299 425
rect 1249 375 1257 409
rect 1291 375 1299 409
rect 1081 307 1089 341
rect 1123 323 1131 341
rect 1249 341 1299 375
rect 1333 409 1383 443
rect 1501 443 1509 459
rect 1543 459 1677 477
rect 1543 443 1551 459
rect 1333 375 1341 409
rect 1375 375 1383 409
rect 1333 357 1383 375
rect 1417 409 1467 425
rect 1417 375 1425 409
rect 1459 375 1467 409
rect 1249 323 1257 341
rect 1123 307 1257 323
rect 1291 323 1299 341
rect 1417 341 1467 375
rect 1501 409 1551 443
rect 1669 443 1677 459
rect 1711 443 1719 477
rect 1501 375 1509 409
rect 1543 375 1551 409
rect 1501 357 1551 375
rect 1585 409 1635 425
rect 1585 375 1593 409
rect 1627 375 1635 409
rect 1417 323 1425 341
rect 1291 307 1425 323
rect 1459 323 1467 341
rect 1585 341 1635 375
rect 1669 409 1719 443
rect 1669 375 1677 409
rect 1711 375 1719 409
rect 1669 357 1719 375
rect 1585 323 1593 341
rect 1459 307 1593 323
rect 1627 323 1635 341
rect 1627 307 1731 323
rect 149 257 183 291
rect 1081 289 1731 307
rect 17 249 115 257
rect 17 215 55 249
rect 89 215 115 249
rect 17 213 115 215
rect 149 249 1000 257
rect 149 215 397 249
rect 431 215 465 249
rect 499 215 533 249
rect 567 215 601 249
rect 635 215 669 249
rect 703 215 737 249
rect 771 215 805 249
rect 839 215 873 249
rect 907 215 941 249
rect 975 215 1000 249
rect 1054 249 1602 255
rect 1054 215 1072 249
rect 1106 215 1140 249
rect 1174 215 1208 249
rect 1242 215 1276 249
rect 1310 215 1344 249
rect 1378 215 1412 249
rect 1446 215 1480 249
rect 1514 215 1548 249
rect 1582 215 1602 249
rect 149 213 231 215
rect 17 51 53 213
rect 87 163 131 179
rect 87 129 97 163
rect 87 95 131 129
rect 87 61 97 95
rect 87 17 131 61
rect 165 163 231 213
rect 1636 181 1731 289
rect 165 129 181 163
rect 215 129 231 163
rect 165 95 231 129
rect 165 61 181 95
rect 215 61 231 95
rect 165 51 231 61
rect 265 163 367 181
rect 265 17 367 61
rect 401 163 1731 181
rect 401 129 417 163
rect 451 145 585 163
rect 451 129 467 145
rect 401 95 467 129
rect 569 129 585 145
rect 619 145 753 163
rect 619 129 635 145
rect 401 61 417 95
rect 451 61 467 95
rect 401 51 467 61
rect 501 95 535 111
rect 501 17 535 61
rect 569 95 635 129
rect 737 129 753 145
rect 787 145 921 163
rect 787 129 803 145
rect 569 61 585 95
rect 619 61 635 95
rect 569 51 635 61
rect 669 95 703 111
rect 669 17 703 61
rect 737 95 803 129
rect 905 129 921 145
rect 955 145 1089 163
rect 955 129 971 145
rect 737 61 753 95
rect 787 61 803 95
rect 737 51 803 61
rect 837 95 871 111
rect 837 17 871 61
rect 905 95 971 129
rect 1073 129 1089 145
rect 1123 145 1257 163
rect 1123 129 1139 145
rect 905 61 921 95
rect 955 61 971 95
rect 905 51 971 61
rect 1005 95 1039 111
rect 1005 17 1039 61
rect 1073 95 1139 129
rect 1241 129 1257 145
rect 1291 145 1425 163
rect 1291 129 1307 145
rect 1073 61 1089 95
rect 1123 61 1139 95
rect 1073 51 1139 61
rect 1173 95 1207 111
rect 1173 17 1207 61
rect 1241 95 1307 129
rect 1409 129 1425 145
rect 1459 145 1593 163
rect 1459 129 1475 145
rect 1241 61 1257 95
rect 1291 61 1307 95
rect 1241 51 1307 61
rect 1341 95 1375 111
rect 1341 17 1375 61
rect 1409 95 1475 129
rect 1577 129 1593 145
rect 1627 145 1731 163
rect 1627 129 1643 145
rect 1409 61 1425 95
rect 1459 61 1475 95
rect 1409 51 1475 61
rect 1509 95 1543 111
rect 1509 17 1543 61
rect 1577 95 1643 129
rect 1577 61 1593 95
rect 1627 61 1643 95
rect 1577 51 1643 61
rect 1677 95 1731 111
rect 1711 61 1731 95
rect 1677 17 1731 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel locali s 37 221 71 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 1670 289 1704 323 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel locali s 1133 221 1167 255 0 FreeSans 400 0 0 0 SLEEP
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 lpflow_isobufsrc_8
rlabel metal1 s 0 -48 1748 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1748 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_END 2398866
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2385564
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 43.700 0.000 
<< end >>
