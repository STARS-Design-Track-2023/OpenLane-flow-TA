magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -66 377 2370 897
<< pwell >>
rect 1865 217 2298 283
rect 8 43 2298 217
rect -26 -43 2330 43
<< locali >>
rect 117 401 359 555
rect 408 437 474 652
rect 117 367 554 401
rect 520 339 554 367
rect 520 289 597 339
rect 703 305 772 499
rect 874 229 933 499
rect 2212 103 2280 751
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2304 831
rect 112 735 302 741
rect 112 701 118 735
rect 152 701 190 735
rect 224 701 262 735
rect 296 701 302 735
rect 26 269 76 679
rect 112 599 302 701
rect 515 569 565 745
rect 673 735 863 745
rect 673 701 679 735
rect 713 701 751 735
rect 785 701 823 735
rect 857 701 863 735
rect 673 605 863 701
rect 899 727 1073 761
rect 899 569 933 727
rect 515 535 933 569
rect 590 381 667 499
rect 393 269 459 331
rect 26 253 459 269
rect 633 253 667 381
rect 806 269 840 535
rect 26 235 667 253
rect 26 99 96 235
rect 393 219 667 235
rect 703 235 840 269
rect 132 113 322 199
rect 703 183 737 235
rect 969 269 1003 691
rect 1039 481 1073 727
rect 1109 735 1143 741
rect 1109 517 1143 701
rect 1179 719 1450 753
rect 1179 481 1213 719
rect 1039 447 1213 481
rect 1249 517 1315 683
rect 1351 585 1450 719
rect 1540 585 1606 751
rect 1737 735 1927 741
rect 1737 701 1743 735
rect 1777 701 1815 735
rect 1849 701 1887 735
rect 1921 701 1927 735
rect 1737 601 1927 701
rect 1979 735 2169 751
rect 1979 701 1985 735
rect 2019 701 2057 735
rect 2091 701 2129 735
rect 2163 701 2169 735
rect 1118 269 1184 369
rect 969 235 1184 269
rect 969 195 1003 235
rect 132 79 138 113
rect 172 79 210 113
rect 244 79 282 113
rect 316 79 322 113
rect 484 149 737 183
rect 484 99 550 149
rect 773 113 891 195
rect 132 73 322 79
rect 773 79 779 113
rect 813 79 851 113
rect 885 79 891 113
rect 939 103 1005 195
rect 1041 113 1159 199
rect 1249 195 1283 517
rect 1351 195 1385 585
rect 1572 565 1606 585
rect 1572 531 1784 565
rect 1568 443 1714 495
rect 1568 351 1602 443
rect 1750 401 1784 531
rect 1877 471 1943 535
rect 1979 507 2169 701
rect 1877 437 2110 471
rect 773 73 891 79
rect 1041 79 1047 113
rect 1081 79 1119 113
rect 1153 79 1159 113
rect 1041 73 1159 79
rect 1209 87 1283 195
rect 1319 123 1385 195
rect 1421 317 1602 351
rect 1638 367 2040 401
rect 1421 87 1455 317
rect 1638 249 1672 367
rect 1974 351 2040 367
rect 1491 215 1672 249
rect 1708 315 1774 331
rect 2076 315 2110 437
rect 1708 281 2110 315
rect 1708 215 1774 281
rect 1491 99 1541 215
rect 1649 113 1839 179
rect 1883 169 1949 281
rect 1209 53 1455 87
rect 1649 79 1655 113
rect 1689 79 1727 113
rect 1761 79 1799 113
rect 1833 79 1839 113
rect 1649 73 1839 79
rect 1985 113 2175 245
rect 1985 79 1991 113
rect 2025 79 2063 113
rect 2097 79 2135 113
rect 2169 79 2175 113
rect 1985 73 2175 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 118 701 152 735
rect 190 701 224 735
rect 262 701 296 735
rect 679 701 713 735
rect 751 701 785 735
rect 823 701 857 735
rect 1109 701 1143 735
rect 1743 701 1777 735
rect 1815 701 1849 735
rect 1887 701 1921 735
rect 1985 701 2019 735
rect 2057 701 2091 735
rect 2129 701 2163 735
rect 138 79 172 113
rect 210 79 244 113
rect 282 79 316 113
rect 779 79 813 113
rect 851 79 885 113
rect 1047 79 1081 113
rect 1119 79 1153 113
rect 1655 79 1689 113
rect 1727 79 1761 113
rect 1799 79 1833 113
rect 1991 79 2025 113
rect 2063 79 2097 113
rect 2135 79 2169 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 831 2304 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2304 831
rect 0 791 2304 797
rect 0 735 2304 763
rect 0 701 118 735
rect 152 701 190 735
rect 224 701 262 735
rect 296 701 679 735
rect 713 701 751 735
rect 785 701 823 735
rect 857 701 1109 735
rect 1143 701 1743 735
rect 1777 701 1815 735
rect 1849 701 1887 735
rect 1921 701 1985 735
rect 2019 701 2057 735
rect 2091 701 2129 735
rect 2163 701 2304 735
rect 0 689 2304 701
rect 0 113 2304 125
rect 0 79 138 113
rect 172 79 210 113
rect 244 79 282 113
rect 316 79 779 113
rect 813 79 851 113
rect 885 79 1047 113
rect 1081 79 1119 113
rect 1153 79 1655 113
rect 1689 79 1727 113
rect 1761 79 1799 113
rect 1833 79 1991 113
rect 2025 79 2063 113
rect 2097 79 2135 113
rect 2169 79 2304 113
rect 0 51 2304 79
rect 0 17 2304 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -23 2304 -17
<< labels >>
rlabel locali s 408 437 474 652 6 D
port 1 nsew signal input
rlabel locali s 874 229 933 499 6 GATE
port 2 nsew clock input
rlabel locali s 703 305 772 499 6 SCD
port 3 nsew signal input
rlabel locali s 520 289 597 339 6 SCE
port 4 nsew signal input
rlabel locali s 520 339 554 367 6 SCE
port 4 nsew signal input
rlabel locali s 117 367 554 401 6 SCE
port 4 nsew signal input
rlabel locali s 117 401 359 555 6 SCE
port 4 nsew signal input
rlabel metal1 s 0 51 2304 125 6 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 -23 2304 23 8 VNB
port 6 nsew ground bidirectional
rlabel pwell s -26 -43 2330 43 8 VNB
port 6 nsew ground bidirectional
rlabel pwell s 8 43 2298 217 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1865 217 2298 283 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 791 2304 837 6 VPB
port 7 nsew power bidirectional
rlabel nwell s -66 377 2370 897 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 689 2304 763 6 VPWR
port 8 nsew power bidirectional
rlabel locali s 2212 103 2280 751 6 Q
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2304 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 719052
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 695106
<< end >>
