magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< dnwell >>
rect 626 14736 14336 36182
<< nwell >>
rect 517 35918 14447 36293
rect 517 15000 832 35918
rect 1593 28312 13423 28975
rect 1593 27622 2336 28312
rect 12680 27622 13423 28312
rect 1593 26878 13423 27622
rect 14072 15000 14447 35918
rect 517 14625 14447 15000
<< pwell >>
rect 219 36363 14750 36600
rect 219 14554 456 36363
rect 1093 34577 13913 34747
rect 1093 15345 1263 34577
rect 13743 15345 13913 34577
rect 1093 15175 13913 15345
rect 14513 14554 14750 36363
rect 219 14317 14750 14554
<< mvpsubdiff >>
rect 245 36497 14724 36574
rect 245 36463 455 36497
rect 489 36463 523 36497
rect 557 36463 591 36497
rect 625 36463 659 36497
rect 693 36463 727 36497
rect 761 36463 795 36497
rect 829 36463 863 36497
rect 897 36463 931 36497
rect 965 36463 999 36497
rect 1033 36463 1067 36497
rect 1101 36463 1135 36497
rect 1169 36463 1203 36497
rect 1237 36463 1271 36497
rect 1305 36463 1339 36497
rect 1373 36463 1407 36497
rect 1441 36463 1475 36497
rect 1509 36463 1543 36497
rect 1577 36463 1611 36497
rect 1645 36463 1679 36497
rect 1713 36463 1747 36497
rect 1781 36463 1815 36497
rect 1849 36463 1883 36497
rect 1917 36463 1951 36497
rect 1985 36463 2019 36497
rect 2053 36463 2087 36497
rect 2121 36463 2155 36497
rect 2189 36463 2223 36497
rect 2257 36463 2291 36497
rect 2325 36463 2359 36497
rect 2393 36463 2427 36497
rect 2461 36463 2495 36497
rect 2529 36463 2563 36497
rect 2597 36463 2631 36497
rect 2665 36463 2699 36497
rect 2733 36463 2767 36497
rect 2801 36463 2835 36497
rect 2869 36463 2903 36497
rect 2937 36463 2971 36497
rect 3005 36463 3039 36497
rect 3073 36463 3107 36497
rect 3141 36463 3175 36497
rect 3209 36463 3243 36497
rect 3277 36463 3311 36497
rect 3345 36463 3379 36497
rect 3413 36463 3447 36497
rect 3481 36463 3515 36497
rect 3549 36463 3583 36497
rect 3617 36463 3651 36497
rect 3685 36463 3719 36497
rect 3753 36463 3787 36497
rect 3821 36463 3855 36497
rect 3889 36463 3923 36497
rect 3957 36463 3991 36497
rect 4025 36463 4059 36497
rect 4093 36463 4127 36497
rect 4161 36463 4195 36497
rect 4229 36463 4263 36497
rect 4297 36463 4331 36497
rect 4365 36463 4399 36497
rect 4433 36463 4467 36497
rect 4501 36463 4535 36497
rect 4569 36463 4603 36497
rect 4637 36463 4671 36497
rect 4705 36463 4739 36497
rect 4773 36463 4807 36497
rect 4841 36463 4875 36497
rect 4909 36463 4943 36497
rect 4977 36463 5011 36497
rect 5045 36463 5079 36497
rect 5113 36463 5147 36497
rect 5181 36463 5215 36497
rect 5249 36463 5283 36497
rect 5317 36463 5351 36497
rect 5385 36463 5419 36497
rect 5453 36463 5487 36497
rect 5521 36463 5555 36497
rect 5589 36463 5623 36497
rect 5657 36463 5691 36497
rect 5725 36463 5759 36497
rect 5793 36463 5827 36497
rect 5861 36463 5895 36497
rect 5929 36463 5963 36497
rect 5997 36463 6031 36497
rect 6065 36463 6099 36497
rect 6133 36463 6167 36497
rect 6201 36463 6235 36497
rect 6269 36463 6303 36497
rect 6337 36463 6371 36497
rect 6405 36463 6439 36497
rect 6473 36463 6507 36497
rect 6541 36463 6575 36497
rect 6609 36463 6643 36497
rect 6677 36463 6711 36497
rect 6745 36463 6779 36497
rect 6813 36463 6847 36497
rect 6881 36463 6915 36497
rect 6949 36463 6983 36497
rect 7017 36463 7051 36497
rect 7085 36463 7119 36497
rect 7153 36463 7187 36497
rect 7221 36463 7255 36497
rect 7289 36463 7323 36497
rect 7357 36463 7391 36497
rect 7425 36463 7459 36497
rect 7493 36463 7527 36497
rect 7561 36463 7595 36497
rect 7629 36463 7663 36497
rect 7697 36463 7731 36497
rect 7765 36463 7799 36497
rect 7833 36463 7867 36497
rect 7901 36463 7935 36497
rect 7969 36463 8003 36497
rect 8037 36463 8071 36497
rect 8105 36463 8139 36497
rect 8173 36463 8207 36497
rect 8241 36463 8275 36497
rect 8309 36463 8343 36497
rect 8377 36463 8411 36497
rect 8445 36463 8479 36497
rect 8513 36463 8547 36497
rect 8581 36463 8615 36497
rect 8649 36463 8683 36497
rect 8717 36463 8751 36497
rect 8785 36463 8819 36497
rect 8853 36463 8887 36497
rect 8921 36463 8955 36497
rect 8989 36463 9023 36497
rect 9057 36463 9091 36497
rect 9125 36463 9159 36497
rect 9193 36463 9227 36497
rect 9261 36463 9295 36497
rect 9329 36463 9363 36497
rect 9397 36463 9431 36497
rect 9465 36463 9499 36497
rect 9533 36463 9567 36497
rect 9601 36463 9635 36497
rect 9669 36463 9703 36497
rect 9737 36463 9771 36497
rect 9805 36463 9839 36497
rect 9873 36463 9907 36497
rect 9941 36463 9975 36497
rect 10009 36463 10043 36497
rect 10077 36463 10111 36497
rect 10145 36463 10179 36497
rect 10213 36463 10247 36497
rect 10281 36463 10315 36497
rect 10349 36463 10383 36497
rect 10417 36463 10451 36497
rect 10485 36463 10519 36497
rect 10553 36463 10587 36497
rect 10621 36463 10655 36497
rect 10689 36463 10723 36497
rect 10757 36463 10791 36497
rect 10825 36463 10859 36497
rect 10893 36463 10927 36497
rect 10961 36463 10995 36497
rect 11029 36463 11063 36497
rect 11097 36463 11131 36497
rect 11165 36463 11199 36497
rect 11233 36463 11267 36497
rect 11301 36463 11335 36497
rect 11369 36463 11403 36497
rect 11437 36463 11471 36497
rect 11505 36463 11539 36497
rect 11573 36463 11607 36497
rect 11641 36463 11675 36497
rect 11709 36463 11743 36497
rect 11777 36463 11811 36497
rect 11845 36463 11879 36497
rect 11913 36463 11947 36497
rect 11981 36463 12015 36497
rect 12049 36463 12083 36497
rect 12117 36463 12151 36497
rect 12185 36463 12219 36497
rect 12253 36463 12287 36497
rect 12321 36463 12355 36497
rect 12389 36463 12423 36497
rect 12457 36463 12491 36497
rect 12525 36463 12559 36497
rect 12593 36463 12627 36497
rect 12661 36463 12695 36497
rect 12729 36463 12763 36497
rect 12797 36463 12831 36497
rect 12865 36463 12899 36497
rect 12933 36463 12967 36497
rect 13001 36463 13035 36497
rect 13069 36463 13103 36497
rect 13137 36463 13171 36497
rect 13205 36463 13239 36497
rect 13273 36463 13307 36497
rect 13341 36463 13375 36497
rect 13409 36463 13443 36497
rect 13477 36463 13511 36497
rect 13545 36463 13579 36497
rect 13613 36463 13647 36497
rect 13681 36463 13715 36497
rect 13749 36463 13783 36497
rect 13817 36463 13851 36497
rect 13885 36463 13919 36497
rect 13953 36463 13987 36497
rect 14021 36463 14055 36497
rect 14089 36463 14123 36497
rect 14157 36463 14191 36497
rect 14225 36463 14259 36497
rect 14293 36463 14327 36497
rect 14361 36463 14395 36497
rect 14429 36463 14463 36497
rect 14497 36463 14724 36497
rect 245 36389 14724 36463
rect 245 36356 430 36389
rect 245 36322 312 36356
rect 346 36322 430 36356
rect 245 36288 430 36322
rect 245 36254 312 36288
rect 346 36254 430 36288
rect 245 36220 430 36254
rect 14539 36362 14724 36389
rect 14539 36328 14607 36362
rect 14641 36328 14724 36362
rect 14539 36294 14724 36328
rect 14539 36260 14607 36294
rect 14641 36260 14724 36294
rect 245 36186 312 36220
rect 346 36186 430 36220
rect 245 36152 430 36186
rect 245 36118 312 36152
rect 346 36118 430 36152
rect 245 36084 430 36118
rect 245 36050 312 36084
rect 346 36050 430 36084
rect 245 36016 430 36050
rect 245 35982 312 36016
rect 346 35982 430 36016
rect 245 35948 430 35982
rect 245 35914 312 35948
rect 346 35914 430 35948
rect 245 35880 430 35914
rect 245 35846 312 35880
rect 346 35846 430 35880
rect 245 35812 430 35846
rect 245 35778 312 35812
rect 346 35778 430 35812
rect 245 35744 430 35778
rect 245 35710 312 35744
rect 346 35710 430 35744
rect 245 35676 430 35710
rect 245 35642 312 35676
rect 346 35642 430 35676
rect 245 35608 430 35642
rect 245 35574 312 35608
rect 346 35574 430 35608
rect 245 35540 430 35574
rect 245 35506 312 35540
rect 346 35506 430 35540
rect 245 35472 430 35506
rect 245 35438 312 35472
rect 346 35438 430 35472
rect 245 35404 430 35438
rect 245 35370 312 35404
rect 346 35370 430 35404
rect 245 35336 430 35370
rect 245 35302 312 35336
rect 346 35302 430 35336
rect 245 35268 430 35302
rect 245 35234 312 35268
rect 346 35234 430 35268
rect 245 35200 430 35234
rect 245 35166 312 35200
rect 346 35166 430 35200
rect 245 35132 430 35166
rect 245 35098 312 35132
rect 346 35098 430 35132
rect 245 35064 430 35098
rect 245 35030 312 35064
rect 346 35030 430 35064
rect 245 34996 430 35030
rect 245 34962 312 34996
rect 346 34962 430 34996
rect 245 34928 430 34962
rect 245 34894 312 34928
rect 346 34894 430 34928
rect 245 34860 430 34894
rect 245 34826 312 34860
rect 346 34826 430 34860
rect 245 34792 430 34826
rect 245 34758 312 34792
rect 346 34758 430 34792
rect 245 34724 430 34758
rect 245 34690 312 34724
rect 346 34690 430 34724
rect 245 34656 430 34690
rect 245 34622 312 34656
rect 346 34622 430 34656
rect 245 34588 430 34622
rect 245 34554 312 34588
rect 346 34554 430 34588
rect 245 34520 430 34554
rect 245 34486 312 34520
rect 346 34486 430 34520
rect 245 34452 430 34486
rect 245 34418 312 34452
rect 346 34418 430 34452
rect 245 34384 430 34418
rect 245 34350 312 34384
rect 346 34350 430 34384
rect 245 34316 430 34350
rect 245 34282 312 34316
rect 346 34282 430 34316
rect 245 34248 430 34282
rect 245 34214 312 34248
rect 346 34214 430 34248
rect 245 34180 430 34214
rect 245 34146 312 34180
rect 346 34146 430 34180
rect 245 34112 430 34146
rect 245 34078 312 34112
rect 346 34078 430 34112
rect 245 34044 430 34078
rect 245 34010 312 34044
rect 346 34010 430 34044
rect 245 33976 430 34010
rect 245 33942 312 33976
rect 346 33942 430 33976
rect 245 33908 430 33942
rect 245 33874 312 33908
rect 346 33874 430 33908
rect 245 33840 430 33874
rect 245 33806 312 33840
rect 346 33806 430 33840
rect 245 33772 430 33806
rect 245 33738 312 33772
rect 346 33738 430 33772
rect 245 33704 430 33738
rect 245 33670 312 33704
rect 346 33670 430 33704
rect 245 33636 430 33670
rect 245 33602 312 33636
rect 346 33602 430 33636
rect 245 33568 430 33602
rect 245 33534 312 33568
rect 346 33534 430 33568
rect 245 33500 430 33534
rect 245 33466 312 33500
rect 346 33466 430 33500
rect 245 33432 430 33466
rect 245 33398 312 33432
rect 346 33398 430 33432
rect 245 33364 430 33398
rect 245 33330 312 33364
rect 346 33330 430 33364
rect 245 33296 430 33330
rect 245 33262 312 33296
rect 346 33262 430 33296
rect 245 33228 430 33262
rect 245 33194 312 33228
rect 346 33194 430 33228
rect 245 33160 430 33194
rect 245 33126 312 33160
rect 346 33126 430 33160
rect 245 33092 430 33126
rect 245 33058 312 33092
rect 346 33058 430 33092
rect 245 33024 430 33058
rect 245 32990 312 33024
rect 346 32990 430 33024
rect 245 32956 430 32990
rect 245 32922 312 32956
rect 346 32922 430 32956
rect 245 32888 430 32922
rect 245 32854 312 32888
rect 346 32854 430 32888
rect 245 32820 430 32854
rect 245 32786 312 32820
rect 346 32786 430 32820
rect 245 32752 430 32786
rect 245 32718 312 32752
rect 346 32718 430 32752
rect 245 32684 430 32718
rect 245 32650 312 32684
rect 346 32650 430 32684
rect 245 32616 430 32650
rect 245 32582 312 32616
rect 346 32582 430 32616
rect 245 32548 430 32582
rect 245 32514 312 32548
rect 346 32514 430 32548
rect 245 32480 430 32514
rect 245 32446 312 32480
rect 346 32446 430 32480
rect 245 32412 430 32446
rect 245 32378 312 32412
rect 346 32378 430 32412
rect 245 32344 430 32378
rect 245 32310 312 32344
rect 346 32310 430 32344
rect 245 32276 430 32310
rect 245 32242 312 32276
rect 346 32242 430 32276
rect 245 32208 430 32242
rect 245 32174 312 32208
rect 346 32174 430 32208
rect 245 32140 430 32174
rect 245 32106 312 32140
rect 346 32106 430 32140
rect 245 32072 430 32106
rect 245 32038 312 32072
rect 346 32038 430 32072
rect 245 32004 430 32038
rect 245 31970 312 32004
rect 346 31970 430 32004
rect 245 31936 430 31970
rect 245 31902 312 31936
rect 346 31902 430 31936
rect 245 31868 430 31902
rect 245 31834 312 31868
rect 346 31834 430 31868
rect 245 31800 430 31834
rect 245 31766 312 31800
rect 346 31766 430 31800
rect 245 31732 430 31766
rect 245 31698 312 31732
rect 346 31698 430 31732
rect 245 31664 430 31698
rect 245 31630 312 31664
rect 346 31630 430 31664
rect 245 31596 430 31630
rect 245 31562 312 31596
rect 346 31562 430 31596
rect 245 31528 430 31562
rect 245 31494 312 31528
rect 346 31494 430 31528
rect 245 31460 430 31494
rect 245 31426 312 31460
rect 346 31426 430 31460
rect 245 31392 430 31426
rect 245 31358 312 31392
rect 346 31358 430 31392
rect 245 31324 430 31358
rect 245 31290 312 31324
rect 346 31290 430 31324
rect 245 31256 430 31290
rect 245 31222 312 31256
rect 346 31222 430 31256
rect 245 31188 430 31222
rect 245 31154 312 31188
rect 346 31154 430 31188
rect 245 31120 430 31154
rect 245 31086 312 31120
rect 346 31086 430 31120
rect 245 31052 430 31086
rect 245 31018 312 31052
rect 346 31018 430 31052
rect 245 30984 430 31018
rect 245 30950 312 30984
rect 346 30950 430 30984
rect 245 30916 430 30950
rect 245 30882 312 30916
rect 346 30882 430 30916
rect 245 30848 430 30882
rect 245 30814 312 30848
rect 346 30814 430 30848
rect 245 30780 430 30814
rect 245 30746 312 30780
rect 346 30746 430 30780
rect 245 30712 430 30746
rect 245 30678 312 30712
rect 346 30678 430 30712
rect 245 30644 430 30678
rect 245 30610 312 30644
rect 346 30610 430 30644
rect 245 30576 430 30610
rect 245 30542 312 30576
rect 346 30542 430 30576
rect 245 30508 430 30542
rect 245 30474 312 30508
rect 346 30474 430 30508
rect 245 30440 430 30474
rect 245 30406 312 30440
rect 346 30406 430 30440
rect 245 30372 430 30406
rect 245 30338 312 30372
rect 346 30338 430 30372
rect 245 30304 430 30338
rect 245 30270 312 30304
rect 346 30270 430 30304
rect 245 30236 430 30270
rect 245 30202 312 30236
rect 346 30202 430 30236
rect 245 30168 430 30202
rect 245 30134 312 30168
rect 346 30134 430 30168
rect 245 30100 430 30134
rect 245 30066 312 30100
rect 346 30066 430 30100
rect 245 30032 430 30066
rect 245 29998 312 30032
rect 346 29998 430 30032
rect 245 29964 430 29998
rect 245 29930 312 29964
rect 346 29930 430 29964
rect 245 29896 430 29930
rect 245 29862 312 29896
rect 346 29862 430 29896
rect 245 29828 430 29862
rect 245 29794 312 29828
rect 346 29794 430 29828
rect 245 29760 430 29794
rect 245 29726 312 29760
rect 346 29726 430 29760
rect 245 29692 430 29726
rect 245 29658 312 29692
rect 346 29658 430 29692
rect 245 29624 430 29658
rect 245 29590 312 29624
rect 346 29590 430 29624
rect 245 29556 430 29590
rect 245 29522 312 29556
rect 346 29522 430 29556
rect 245 29488 430 29522
rect 245 29454 312 29488
rect 346 29454 430 29488
rect 245 29420 430 29454
rect 245 29386 312 29420
rect 346 29386 430 29420
rect 245 29352 430 29386
rect 245 29318 312 29352
rect 346 29318 430 29352
rect 245 29284 430 29318
rect 245 29250 312 29284
rect 346 29250 430 29284
rect 245 29216 430 29250
rect 245 29182 312 29216
rect 346 29182 430 29216
rect 245 29148 430 29182
rect 245 29114 312 29148
rect 346 29114 430 29148
rect 245 29080 430 29114
rect 245 29046 312 29080
rect 346 29046 430 29080
rect 245 29012 430 29046
rect 245 28978 312 29012
rect 346 28978 430 29012
rect 245 28944 430 28978
rect 245 28910 312 28944
rect 346 28910 430 28944
rect 245 28876 430 28910
rect 245 28842 312 28876
rect 346 28842 430 28876
rect 245 28808 430 28842
rect 245 28774 312 28808
rect 346 28774 430 28808
rect 245 28740 430 28774
rect 245 28706 312 28740
rect 346 28706 430 28740
rect 245 28672 430 28706
rect 245 28638 312 28672
rect 346 28638 430 28672
rect 245 28604 430 28638
rect 245 28570 312 28604
rect 346 28570 430 28604
rect 245 28536 430 28570
rect 245 28502 312 28536
rect 346 28502 430 28536
rect 245 28468 430 28502
rect 245 28434 312 28468
rect 346 28434 430 28468
rect 245 28400 430 28434
rect 245 28366 312 28400
rect 346 28366 430 28400
rect 245 28332 430 28366
rect 245 28298 312 28332
rect 346 28298 430 28332
rect 245 28264 430 28298
rect 245 28230 312 28264
rect 346 28230 430 28264
rect 245 28196 430 28230
rect 245 28162 312 28196
rect 346 28162 430 28196
rect 245 28128 430 28162
rect 245 28094 312 28128
rect 346 28094 430 28128
rect 245 28060 430 28094
rect 245 28026 312 28060
rect 346 28026 430 28060
rect 245 27992 430 28026
rect 245 27958 312 27992
rect 346 27958 430 27992
rect 245 27924 430 27958
rect 245 27890 312 27924
rect 346 27890 430 27924
rect 245 27856 430 27890
rect 245 27822 312 27856
rect 346 27822 430 27856
rect 245 27788 430 27822
rect 245 27754 312 27788
rect 346 27754 430 27788
rect 245 27720 430 27754
rect 245 27686 312 27720
rect 346 27686 430 27720
rect 245 27652 430 27686
rect 245 27618 312 27652
rect 346 27618 430 27652
rect 245 27584 430 27618
rect 245 27550 312 27584
rect 346 27550 430 27584
rect 245 27516 430 27550
rect 245 27482 312 27516
rect 346 27482 430 27516
rect 245 27448 430 27482
rect 245 27414 312 27448
rect 346 27414 430 27448
rect 245 27380 430 27414
rect 245 27346 312 27380
rect 346 27346 430 27380
rect 245 27312 430 27346
rect 245 27278 312 27312
rect 346 27278 430 27312
rect 245 27244 430 27278
rect 245 27210 312 27244
rect 346 27210 430 27244
rect 245 27176 430 27210
rect 245 27142 312 27176
rect 346 27142 430 27176
rect 245 27108 430 27142
rect 245 27074 312 27108
rect 346 27074 430 27108
rect 245 27040 430 27074
rect 245 27006 312 27040
rect 346 27006 430 27040
rect 245 26972 430 27006
rect 245 26938 312 26972
rect 346 26938 430 26972
rect 245 26904 430 26938
rect 245 26870 312 26904
rect 346 26870 430 26904
rect 245 26836 430 26870
rect 245 26802 312 26836
rect 346 26802 430 26836
rect 245 26768 430 26802
rect 245 26734 312 26768
rect 346 26734 430 26768
rect 245 26700 430 26734
rect 245 26666 312 26700
rect 346 26666 430 26700
rect 245 26632 430 26666
rect 245 26598 312 26632
rect 346 26598 430 26632
rect 245 26564 430 26598
rect 245 26530 312 26564
rect 346 26530 430 26564
rect 245 26496 430 26530
rect 245 26462 312 26496
rect 346 26462 430 26496
rect 245 26428 430 26462
rect 245 26394 312 26428
rect 346 26394 430 26428
rect 245 26360 430 26394
rect 245 26326 312 26360
rect 346 26326 430 26360
rect 245 26292 430 26326
rect 245 26258 312 26292
rect 346 26258 430 26292
rect 245 26224 430 26258
rect 245 26190 312 26224
rect 346 26190 430 26224
rect 245 26156 430 26190
rect 245 26122 312 26156
rect 346 26122 430 26156
rect 245 26088 430 26122
rect 245 26054 312 26088
rect 346 26054 430 26088
rect 245 26020 430 26054
rect 245 25986 312 26020
rect 346 25986 430 26020
rect 245 25952 430 25986
rect 245 25918 312 25952
rect 346 25918 430 25952
rect 245 25884 430 25918
rect 245 25850 312 25884
rect 346 25850 430 25884
rect 245 25816 430 25850
rect 245 25782 312 25816
rect 346 25782 430 25816
rect 245 25748 430 25782
rect 245 25714 312 25748
rect 346 25714 430 25748
rect 245 25680 430 25714
rect 245 25646 312 25680
rect 346 25646 430 25680
rect 245 25612 430 25646
rect 245 25578 312 25612
rect 346 25578 430 25612
rect 245 25544 430 25578
rect 245 25510 312 25544
rect 346 25510 430 25544
rect 245 25476 430 25510
rect 245 25442 312 25476
rect 346 25442 430 25476
rect 245 25408 430 25442
rect 245 25374 312 25408
rect 346 25374 430 25408
rect 245 25340 430 25374
rect 245 25306 312 25340
rect 346 25306 430 25340
rect 245 25272 430 25306
rect 245 25238 312 25272
rect 346 25238 430 25272
rect 245 25204 430 25238
rect 245 25170 312 25204
rect 346 25170 430 25204
rect 245 25136 430 25170
rect 245 25102 312 25136
rect 346 25102 430 25136
rect 245 25068 430 25102
rect 245 25034 312 25068
rect 346 25034 430 25068
rect 245 25000 430 25034
rect 245 24966 312 25000
rect 346 24966 430 25000
rect 245 24932 430 24966
rect 245 24898 312 24932
rect 346 24898 430 24932
rect 245 24864 430 24898
rect 245 24830 312 24864
rect 346 24830 430 24864
rect 245 24796 430 24830
rect 245 24762 312 24796
rect 346 24762 430 24796
rect 245 24728 430 24762
rect 245 24694 312 24728
rect 346 24694 430 24728
rect 245 24660 430 24694
rect 245 24626 312 24660
rect 346 24626 430 24660
rect 245 24592 430 24626
rect 245 24558 312 24592
rect 346 24558 430 24592
rect 245 24524 430 24558
rect 245 24490 312 24524
rect 346 24490 430 24524
rect 245 24456 430 24490
rect 245 24422 312 24456
rect 346 24422 430 24456
rect 245 24388 430 24422
rect 245 24354 312 24388
rect 346 24354 430 24388
rect 245 24320 430 24354
rect 245 24286 312 24320
rect 346 24286 430 24320
rect 245 24252 430 24286
rect 245 24218 312 24252
rect 346 24218 430 24252
rect 245 24184 430 24218
rect 245 24150 312 24184
rect 346 24150 430 24184
rect 245 24116 430 24150
rect 245 24082 312 24116
rect 346 24082 430 24116
rect 245 24048 430 24082
rect 245 24014 312 24048
rect 346 24014 430 24048
rect 245 23980 430 24014
rect 245 23946 312 23980
rect 346 23946 430 23980
rect 245 23912 430 23946
rect 245 23878 312 23912
rect 346 23878 430 23912
rect 245 23844 430 23878
rect 245 23810 312 23844
rect 346 23810 430 23844
rect 245 23776 430 23810
rect 245 23742 312 23776
rect 346 23742 430 23776
rect 245 23708 430 23742
rect 245 23674 312 23708
rect 346 23674 430 23708
rect 245 23640 430 23674
rect 245 23606 312 23640
rect 346 23606 430 23640
rect 245 23572 430 23606
rect 245 23538 312 23572
rect 346 23538 430 23572
rect 245 23504 430 23538
rect 245 23470 312 23504
rect 346 23470 430 23504
rect 245 23436 430 23470
rect 245 23402 312 23436
rect 346 23402 430 23436
rect 245 23368 430 23402
rect 245 23334 312 23368
rect 346 23334 430 23368
rect 245 23300 430 23334
rect 245 23266 312 23300
rect 346 23266 430 23300
rect 245 23232 430 23266
rect 245 23198 312 23232
rect 346 23198 430 23232
rect 245 23164 430 23198
rect 245 23130 312 23164
rect 346 23130 430 23164
rect 245 23096 430 23130
rect 245 23062 312 23096
rect 346 23062 430 23096
rect 245 23028 430 23062
rect 245 22994 312 23028
rect 346 22994 430 23028
rect 245 22960 430 22994
rect 245 22926 312 22960
rect 346 22926 430 22960
rect 245 22892 430 22926
rect 245 22858 312 22892
rect 346 22858 430 22892
rect 245 22824 430 22858
rect 245 22790 312 22824
rect 346 22790 430 22824
rect 245 22756 430 22790
rect 245 22722 312 22756
rect 346 22722 430 22756
rect 245 22688 430 22722
rect 245 22654 312 22688
rect 346 22654 430 22688
rect 245 22620 430 22654
rect 245 22586 312 22620
rect 346 22586 430 22620
rect 245 22552 430 22586
rect 245 22518 312 22552
rect 346 22518 430 22552
rect 245 22484 430 22518
rect 245 22450 312 22484
rect 346 22450 430 22484
rect 245 22416 430 22450
rect 245 22382 312 22416
rect 346 22382 430 22416
rect 245 22348 430 22382
rect 245 22314 312 22348
rect 346 22314 430 22348
rect 245 22280 430 22314
rect 245 22246 312 22280
rect 346 22246 430 22280
rect 245 22212 430 22246
rect 245 22178 312 22212
rect 346 22178 430 22212
rect 245 22144 430 22178
rect 245 22110 312 22144
rect 346 22110 430 22144
rect 245 22076 430 22110
rect 245 22042 312 22076
rect 346 22042 430 22076
rect 245 22008 430 22042
rect 245 21974 312 22008
rect 346 21974 430 22008
rect 245 21940 430 21974
rect 245 21906 312 21940
rect 346 21906 430 21940
rect 245 21872 430 21906
rect 245 21838 312 21872
rect 346 21838 430 21872
rect 245 21804 430 21838
rect 245 21770 312 21804
rect 346 21770 430 21804
rect 245 21736 430 21770
rect 245 21702 312 21736
rect 346 21702 430 21736
rect 245 21668 430 21702
rect 245 21634 312 21668
rect 346 21634 430 21668
rect 245 21600 430 21634
rect 245 21566 312 21600
rect 346 21566 430 21600
rect 245 21532 430 21566
rect 245 21498 312 21532
rect 346 21498 430 21532
rect 245 21464 430 21498
rect 245 21430 312 21464
rect 346 21430 430 21464
rect 245 21396 430 21430
rect 245 21362 312 21396
rect 346 21362 430 21396
rect 245 21328 430 21362
rect 245 21294 312 21328
rect 346 21294 430 21328
rect 245 21260 430 21294
rect 245 21226 312 21260
rect 346 21226 430 21260
rect 245 21192 430 21226
rect 245 21158 312 21192
rect 346 21158 430 21192
rect 245 21124 430 21158
rect 245 21090 312 21124
rect 346 21090 430 21124
rect 245 21056 430 21090
rect 245 21022 312 21056
rect 346 21022 430 21056
rect 245 20988 430 21022
rect 245 20954 312 20988
rect 346 20954 430 20988
rect 245 20920 430 20954
rect 245 20886 312 20920
rect 346 20886 430 20920
rect 245 20852 430 20886
rect 245 20818 312 20852
rect 346 20818 430 20852
rect 245 20784 430 20818
rect 245 20750 312 20784
rect 346 20750 430 20784
rect 245 20716 430 20750
rect 245 20682 312 20716
rect 346 20682 430 20716
rect 245 20648 430 20682
rect 245 20614 312 20648
rect 346 20614 430 20648
rect 245 20580 430 20614
rect 245 20546 312 20580
rect 346 20546 430 20580
rect 245 20512 430 20546
rect 245 20478 312 20512
rect 346 20478 430 20512
rect 245 20444 430 20478
rect 245 20410 312 20444
rect 346 20410 430 20444
rect 245 20376 430 20410
rect 245 20342 312 20376
rect 346 20342 430 20376
rect 245 20308 430 20342
rect 245 20274 312 20308
rect 346 20274 430 20308
rect 245 20240 430 20274
rect 245 20206 312 20240
rect 346 20206 430 20240
rect 245 20172 430 20206
rect 245 20138 312 20172
rect 346 20138 430 20172
rect 245 20104 430 20138
rect 245 20070 312 20104
rect 346 20070 430 20104
rect 245 20036 430 20070
rect 245 20002 312 20036
rect 346 20002 430 20036
rect 245 19968 430 20002
rect 245 19934 312 19968
rect 346 19934 430 19968
rect 245 19900 430 19934
rect 245 19866 312 19900
rect 346 19866 430 19900
rect 245 19832 430 19866
rect 245 19798 312 19832
rect 346 19798 430 19832
rect 245 19764 430 19798
rect 245 19730 312 19764
rect 346 19730 430 19764
rect 245 19696 430 19730
rect 245 19662 312 19696
rect 346 19662 430 19696
rect 245 19628 430 19662
rect 245 19594 312 19628
rect 346 19594 430 19628
rect 245 19560 430 19594
rect 245 19526 312 19560
rect 346 19526 430 19560
rect 245 19492 430 19526
rect 245 19458 312 19492
rect 346 19458 430 19492
rect 245 19424 430 19458
rect 245 19390 312 19424
rect 346 19390 430 19424
rect 245 19356 430 19390
rect 245 19322 312 19356
rect 346 19322 430 19356
rect 245 19288 430 19322
rect 245 19254 312 19288
rect 346 19254 430 19288
rect 245 19220 430 19254
rect 245 19186 312 19220
rect 346 19186 430 19220
rect 245 19152 430 19186
rect 245 19118 312 19152
rect 346 19118 430 19152
rect 245 19084 430 19118
rect 245 19050 312 19084
rect 346 19050 430 19084
rect 245 19016 430 19050
rect 245 18982 312 19016
rect 346 18982 430 19016
rect 245 18948 430 18982
rect 245 18914 312 18948
rect 346 18914 430 18948
rect 245 18880 430 18914
rect 245 18846 312 18880
rect 346 18846 430 18880
rect 245 18812 430 18846
rect 245 18778 312 18812
rect 346 18778 430 18812
rect 245 18744 430 18778
rect 245 18710 312 18744
rect 346 18710 430 18744
rect 245 18676 430 18710
rect 245 18642 312 18676
rect 346 18642 430 18676
rect 245 18608 430 18642
rect 245 18574 312 18608
rect 346 18574 430 18608
rect 245 18540 430 18574
rect 245 18506 312 18540
rect 346 18506 430 18540
rect 245 18472 430 18506
rect 245 18438 312 18472
rect 346 18438 430 18472
rect 245 18404 430 18438
rect 245 18370 312 18404
rect 346 18370 430 18404
rect 245 18336 430 18370
rect 245 18302 312 18336
rect 346 18302 430 18336
rect 245 18268 430 18302
rect 245 18234 312 18268
rect 346 18234 430 18268
rect 245 18200 430 18234
rect 245 18166 312 18200
rect 346 18166 430 18200
rect 245 18132 430 18166
rect 245 18098 312 18132
rect 346 18098 430 18132
rect 245 18064 430 18098
rect 245 18030 312 18064
rect 346 18030 430 18064
rect 245 17996 430 18030
rect 245 17962 312 17996
rect 346 17962 430 17996
rect 245 17928 430 17962
rect 245 17894 312 17928
rect 346 17894 430 17928
rect 245 17860 430 17894
rect 245 17826 312 17860
rect 346 17826 430 17860
rect 245 17792 430 17826
rect 245 17758 312 17792
rect 346 17758 430 17792
rect 245 17724 430 17758
rect 245 17690 312 17724
rect 346 17690 430 17724
rect 245 17656 430 17690
rect 245 17622 312 17656
rect 346 17622 430 17656
rect 245 17588 430 17622
rect 245 17554 312 17588
rect 346 17554 430 17588
rect 245 17520 430 17554
rect 245 17486 312 17520
rect 346 17486 430 17520
rect 245 17452 430 17486
rect 245 17418 312 17452
rect 346 17418 430 17452
rect 245 17384 430 17418
rect 245 17350 312 17384
rect 346 17350 430 17384
rect 245 17316 430 17350
rect 245 17282 312 17316
rect 346 17282 430 17316
rect 245 17248 430 17282
rect 245 17214 312 17248
rect 346 17214 430 17248
rect 245 17180 430 17214
rect 245 17146 312 17180
rect 346 17146 430 17180
rect 245 17112 430 17146
rect 245 17078 312 17112
rect 346 17078 430 17112
rect 245 17044 430 17078
rect 245 17010 312 17044
rect 346 17010 430 17044
rect 245 16976 430 17010
rect 245 16942 312 16976
rect 346 16942 430 16976
rect 245 16908 430 16942
rect 245 16874 312 16908
rect 346 16874 430 16908
rect 245 16840 430 16874
rect 245 16806 312 16840
rect 346 16806 430 16840
rect 245 16772 430 16806
rect 245 16738 312 16772
rect 346 16738 430 16772
rect 245 16704 430 16738
rect 245 16670 312 16704
rect 346 16670 430 16704
rect 245 16636 430 16670
rect 245 16602 312 16636
rect 346 16602 430 16636
rect 245 16568 430 16602
rect 245 16534 312 16568
rect 346 16534 430 16568
rect 245 16500 430 16534
rect 245 16466 312 16500
rect 346 16466 430 16500
rect 245 16432 430 16466
rect 245 16398 312 16432
rect 346 16398 430 16432
rect 245 16364 430 16398
rect 245 16330 312 16364
rect 346 16330 430 16364
rect 245 16296 430 16330
rect 245 16262 312 16296
rect 346 16262 430 16296
rect 245 16228 430 16262
rect 245 16194 312 16228
rect 346 16194 430 16228
rect 245 16160 430 16194
rect 245 16126 312 16160
rect 346 16126 430 16160
rect 245 16092 430 16126
rect 245 16058 312 16092
rect 346 16058 430 16092
rect 245 16024 430 16058
rect 245 15990 312 16024
rect 346 15990 430 16024
rect 245 15956 430 15990
rect 245 15922 312 15956
rect 346 15922 430 15956
rect 245 15888 430 15922
rect 245 15854 312 15888
rect 346 15854 430 15888
rect 245 15820 430 15854
rect 245 15786 312 15820
rect 346 15786 430 15820
rect 245 15752 430 15786
rect 245 15718 312 15752
rect 346 15718 430 15752
rect 245 15684 430 15718
rect 245 15650 312 15684
rect 346 15650 430 15684
rect 245 15616 430 15650
rect 245 15582 312 15616
rect 346 15582 430 15616
rect 245 15548 430 15582
rect 245 15514 312 15548
rect 346 15514 430 15548
rect 245 15480 430 15514
rect 245 15446 312 15480
rect 346 15446 430 15480
rect 245 15412 430 15446
rect 245 15378 312 15412
rect 346 15378 430 15412
rect 245 15344 430 15378
rect 245 15310 312 15344
rect 346 15310 430 15344
rect 245 15276 430 15310
rect 245 15242 312 15276
rect 346 15242 430 15276
rect 245 15208 430 15242
rect 245 15174 312 15208
rect 346 15174 430 15208
rect 245 15140 430 15174
rect 245 15106 312 15140
rect 346 15106 430 15140
rect 245 15072 430 15106
rect 245 15038 312 15072
rect 346 15038 430 15072
rect 245 15004 430 15038
rect 245 14970 312 15004
rect 346 14970 430 15004
rect 245 14936 430 14970
rect 245 14902 312 14936
rect 346 14902 430 14936
rect 245 14868 430 14902
rect 245 14834 312 14868
rect 346 14834 430 14868
rect 245 14800 430 14834
rect 245 14766 312 14800
rect 346 14766 430 14800
rect 245 14732 430 14766
rect 245 14698 312 14732
rect 346 14698 430 14732
rect 245 14664 430 14698
rect 1119 34679 13887 34721
rect 1119 34645 1305 34679
rect 1339 34645 1373 34679
rect 1407 34645 1441 34679
rect 1475 34645 1509 34679
rect 1543 34645 1577 34679
rect 1611 34645 1645 34679
rect 1679 34645 1713 34679
rect 1747 34645 1781 34679
rect 1815 34645 1849 34679
rect 1883 34645 1917 34679
rect 1951 34645 1985 34679
rect 2019 34645 2053 34679
rect 2087 34645 2121 34679
rect 2155 34645 2189 34679
rect 2223 34645 2257 34679
rect 2291 34645 2325 34679
rect 2359 34645 2393 34679
rect 2427 34645 2461 34679
rect 2495 34645 2529 34679
rect 2563 34645 2597 34679
rect 2631 34645 2665 34679
rect 2699 34645 2733 34679
rect 2767 34645 2801 34679
rect 2835 34645 2869 34679
rect 2903 34645 2937 34679
rect 2971 34645 3005 34679
rect 3039 34645 3073 34679
rect 3107 34645 3141 34679
rect 3175 34645 3209 34679
rect 3243 34645 3277 34679
rect 3311 34645 3345 34679
rect 3379 34645 3413 34679
rect 3447 34645 3481 34679
rect 3515 34645 3549 34679
rect 3583 34645 3617 34679
rect 3651 34645 3685 34679
rect 3719 34645 3753 34679
rect 3787 34645 3821 34679
rect 3855 34645 3889 34679
rect 3923 34645 3957 34679
rect 3991 34645 4025 34679
rect 4059 34645 4093 34679
rect 4127 34645 4161 34679
rect 4195 34645 4229 34679
rect 4263 34645 4297 34679
rect 4331 34645 4365 34679
rect 4399 34645 4433 34679
rect 4467 34645 4501 34679
rect 4535 34645 4569 34679
rect 4603 34645 4637 34679
rect 4671 34645 4705 34679
rect 4739 34645 4773 34679
rect 4807 34645 4841 34679
rect 4875 34645 4909 34679
rect 4943 34645 4977 34679
rect 5011 34645 5045 34679
rect 5079 34645 5113 34679
rect 5147 34645 5181 34679
rect 5215 34645 5249 34679
rect 5283 34645 5317 34679
rect 5351 34645 5385 34679
rect 5419 34645 5453 34679
rect 5487 34645 5521 34679
rect 5555 34645 5589 34679
rect 5623 34645 5657 34679
rect 5691 34645 5725 34679
rect 5759 34645 5793 34679
rect 5827 34645 5861 34679
rect 5895 34645 5929 34679
rect 5963 34645 5997 34679
rect 6031 34645 6065 34679
rect 6099 34645 6133 34679
rect 6167 34645 6201 34679
rect 6235 34645 6269 34679
rect 6303 34645 6337 34679
rect 6371 34645 6405 34679
rect 6439 34645 6473 34679
rect 6507 34645 6541 34679
rect 6575 34645 6609 34679
rect 6643 34645 6677 34679
rect 6711 34645 6745 34679
rect 6779 34645 6813 34679
rect 6847 34645 6881 34679
rect 6915 34645 6949 34679
rect 6983 34645 7017 34679
rect 7051 34645 7085 34679
rect 7119 34645 7153 34679
rect 7187 34645 7221 34679
rect 7255 34645 7289 34679
rect 7323 34645 7357 34679
rect 7391 34645 7425 34679
rect 7459 34645 7493 34679
rect 7527 34645 7561 34679
rect 7595 34645 7629 34679
rect 7663 34645 7697 34679
rect 7731 34645 7765 34679
rect 7799 34645 7833 34679
rect 7867 34645 7901 34679
rect 7935 34645 7969 34679
rect 8003 34645 8037 34679
rect 8071 34645 8105 34679
rect 8139 34645 8173 34679
rect 8207 34645 8241 34679
rect 8275 34645 8309 34679
rect 8343 34645 8377 34679
rect 8411 34645 8445 34679
rect 8479 34645 8513 34679
rect 8547 34645 8581 34679
rect 8615 34645 8649 34679
rect 8683 34645 8717 34679
rect 8751 34645 8785 34679
rect 8819 34645 8853 34679
rect 8887 34645 8921 34679
rect 8955 34645 8989 34679
rect 9023 34645 9057 34679
rect 9091 34645 9125 34679
rect 9159 34645 9193 34679
rect 9227 34645 9261 34679
rect 9295 34645 9329 34679
rect 9363 34645 9397 34679
rect 9431 34645 9465 34679
rect 9499 34645 9533 34679
rect 9567 34645 9601 34679
rect 9635 34645 9669 34679
rect 9703 34645 9737 34679
rect 9771 34645 9805 34679
rect 9839 34645 9873 34679
rect 9907 34645 9941 34679
rect 9975 34645 10009 34679
rect 10043 34645 10077 34679
rect 10111 34645 10145 34679
rect 10179 34645 10213 34679
rect 10247 34645 10281 34679
rect 10315 34645 10349 34679
rect 10383 34645 10417 34679
rect 10451 34645 10485 34679
rect 10519 34645 10553 34679
rect 10587 34645 10621 34679
rect 10655 34645 10689 34679
rect 10723 34645 10757 34679
rect 10791 34645 10825 34679
rect 10859 34645 10893 34679
rect 10927 34645 10961 34679
rect 10995 34645 11029 34679
rect 11063 34645 11097 34679
rect 11131 34645 11165 34679
rect 11199 34645 11233 34679
rect 11267 34645 11301 34679
rect 11335 34645 11369 34679
rect 11403 34645 11437 34679
rect 11471 34645 11505 34679
rect 11539 34645 11573 34679
rect 11607 34645 11641 34679
rect 11675 34645 11709 34679
rect 11743 34645 11777 34679
rect 11811 34645 11845 34679
rect 11879 34645 11913 34679
rect 11947 34645 11981 34679
rect 12015 34645 12049 34679
rect 12083 34645 12117 34679
rect 12151 34645 12185 34679
rect 12219 34645 12253 34679
rect 12287 34645 12321 34679
rect 12355 34645 12389 34679
rect 12423 34645 12457 34679
rect 12491 34645 12525 34679
rect 12559 34645 12593 34679
rect 12627 34645 12661 34679
rect 12695 34645 12729 34679
rect 12763 34645 12797 34679
rect 12831 34645 12865 34679
rect 12899 34645 12933 34679
rect 12967 34645 13001 34679
rect 13035 34645 13069 34679
rect 13103 34645 13137 34679
rect 13171 34645 13205 34679
rect 13239 34645 13273 34679
rect 13307 34645 13341 34679
rect 13375 34645 13409 34679
rect 13443 34645 13477 34679
rect 13511 34645 13545 34679
rect 13579 34645 13613 34679
rect 13647 34645 13681 34679
rect 13715 34645 13887 34679
rect 1119 34603 13887 34645
rect 1119 34462 1237 34603
rect 1119 34428 1161 34462
rect 1195 34428 1237 34462
rect 1119 34394 1237 34428
rect 1119 34360 1161 34394
rect 1195 34360 1237 34394
rect 1119 34326 1237 34360
rect 1119 34292 1161 34326
rect 1195 34292 1237 34326
rect 1119 34258 1237 34292
rect 1119 34224 1161 34258
rect 1195 34224 1237 34258
rect 1119 34190 1237 34224
rect 1119 34156 1161 34190
rect 1195 34156 1237 34190
rect 1119 34122 1237 34156
rect 1119 34088 1161 34122
rect 1195 34088 1237 34122
rect 1119 34054 1237 34088
rect 1119 34020 1161 34054
rect 1195 34020 1237 34054
rect 1119 33986 1237 34020
rect 1119 33952 1161 33986
rect 1195 33952 1237 33986
rect 1119 33918 1237 33952
rect 1119 33884 1161 33918
rect 1195 33884 1237 33918
rect 1119 33850 1237 33884
rect 1119 33816 1161 33850
rect 1195 33816 1237 33850
rect 1119 33782 1237 33816
rect 1119 33748 1161 33782
rect 1195 33748 1237 33782
rect 1119 33714 1237 33748
rect 1119 33680 1161 33714
rect 1195 33680 1237 33714
rect 1119 33646 1237 33680
rect 1119 33612 1161 33646
rect 1195 33612 1237 33646
rect 1119 33578 1237 33612
rect 1119 33544 1161 33578
rect 1195 33544 1237 33578
rect 1119 33510 1237 33544
rect 1119 33476 1161 33510
rect 1195 33476 1237 33510
rect 1119 33442 1237 33476
rect 1119 33408 1161 33442
rect 1195 33408 1237 33442
rect 1119 33374 1237 33408
rect 1119 33340 1161 33374
rect 1195 33340 1237 33374
rect 1119 33306 1237 33340
rect 1119 33272 1161 33306
rect 1195 33272 1237 33306
rect 1119 33238 1237 33272
rect 1119 33204 1161 33238
rect 1195 33204 1237 33238
rect 1119 33170 1237 33204
rect 1119 33136 1161 33170
rect 1195 33136 1237 33170
rect 1119 33102 1237 33136
rect 1119 33068 1161 33102
rect 1195 33068 1237 33102
rect 1119 33034 1237 33068
rect 1119 33000 1161 33034
rect 1195 33000 1237 33034
rect 1119 32966 1237 33000
rect 1119 32932 1161 32966
rect 1195 32932 1237 32966
rect 1119 32898 1237 32932
rect 1119 32864 1161 32898
rect 1195 32864 1237 32898
rect 1119 32830 1237 32864
rect 1119 32796 1161 32830
rect 1195 32796 1237 32830
rect 1119 32762 1237 32796
rect 1119 32728 1161 32762
rect 1195 32728 1237 32762
rect 1119 32694 1237 32728
rect 1119 32660 1161 32694
rect 1195 32660 1237 32694
rect 1119 32626 1237 32660
rect 1119 32592 1161 32626
rect 1195 32592 1237 32626
rect 1119 32558 1237 32592
rect 1119 32524 1161 32558
rect 1195 32524 1237 32558
rect 1119 32490 1237 32524
rect 1119 32456 1161 32490
rect 1195 32456 1237 32490
rect 1119 32422 1237 32456
rect 1119 32388 1161 32422
rect 1195 32388 1237 32422
rect 1119 32354 1237 32388
rect 1119 32320 1161 32354
rect 1195 32320 1237 32354
rect 1119 32286 1237 32320
rect 1119 32252 1161 32286
rect 1195 32252 1237 32286
rect 1119 32218 1237 32252
rect 1119 32184 1161 32218
rect 1195 32184 1237 32218
rect 1119 32150 1237 32184
rect 1119 32116 1161 32150
rect 1195 32116 1237 32150
rect 1119 32082 1237 32116
rect 1119 32048 1161 32082
rect 1195 32048 1237 32082
rect 1119 32014 1237 32048
rect 1119 31980 1161 32014
rect 1195 31980 1237 32014
rect 1119 31946 1237 31980
rect 1119 31912 1161 31946
rect 1195 31912 1237 31946
rect 1119 31878 1237 31912
rect 1119 31844 1161 31878
rect 1195 31844 1237 31878
rect 1119 31810 1237 31844
rect 1119 31776 1161 31810
rect 1195 31776 1237 31810
rect 1119 31742 1237 31776
rect 1119 31708 1161 31742
rect 1195 31708 1237 31742
rect 1119 31674 1237 31708
rect 1119 31640 1161 31674
rect 1195 31640 1237 31674
rect 1119 31606 1237 31640
rect 1119 31572 1161 31606
rect 1195 31572 1237 31606
rect 1119 31538 1237 31572
rect 1119 31504 1161 31538
rect 1195 31504 1237 31538
rect 1119 31470 1237 31504
rect 1119 31436 1161 31470
rect 1195 31436 1237 31470
rect 1119 31402 1237 31436
rect 1119 31368 1161 31402
rect 1195 31368 1237 31402
rect 1119 31334 1237 31368
rect 1119 31300 1161 31334
rect 1195 31300 1237 31334
rect 1119 31266 1237 31300
rect 1119 31232 1161 31266
rect 1195 31232 1237 31266
rect 1119 31198 1237 31232
rect 1119 31164 1161 31198
rect 1195 31164 1237 31198
rect 1119 31130 1237 31164
rect 1119 31096 1161 31130
rect 1195 31096 1237 31130
rect 1119 31062 1237 31096
rect 1119 31028 1161 31062
rect 1195 31028 1237 31062
rect 1119 30994 1237 31028
rect 1119 30960 1161 30994
rect 1195 30960 1237 30994
rect 1119 30926 1237 30960
rect 1119 30892 1161 30926
rect 1195 30892 1237 30926
rect 1119 30858 1237 30892
rect 1119 30824 1161 30858
rect 1195 30824 1237 30858
rect 1119 30790 1237 30824
rect 1119 30756 1161 30790
rect 1195 30756 1237 30790
rect 1119 30722 1237 30756
rect 1119 30688 1161 30722
rect 1195 30688 1237 30722
rect 1119 30654 1237 30688
rect 1119 30620 1161 30654
rect 1195 30620 1237 30654
rect 1119 30586 1237 30620
rect 1119 30552 1161 30586
rect 1195 30552 1237 30586
rect 1119 30518 1237 30552
rect 1119 30484 1161 30518
rect 1195 30484 1237 30518
rect 1119 30450 1237 30484
rect 1119 30416 1161 30450
rect 1195 30416 1237 30450
rect 1119 30382 1237 30416
rect 1119 30348 1161 30382
rect 1195 30348 1237 30382
rect 1119 30314 1237 30348
rect 1119 30280 1161 30314
rect 1195 30280 1237 30314
rect 1119 30246 1237 30280
rect 1119 30212 1161 30246
rect 1195 30212 1237 30246
rect 1119 30178 1237 30212
rect 1119 30144 1161 30178
rect 1195 30144 1237 30178
rect 1119 30110 1237 30144
rect 1119 30076 1161 30110
rect 1195 30076 1237 30110
rect 1119 30042 1237 30076
rect 1119 30008 1161 30042
rect 1195 30008 1237 30042
rect 1119 29974 1237 30008
rect 1119 29940 1161 29974
rect 1195 29940 1237 29974
rect 1119 29906 1237 29940
rect 1119 29872 1161 29906
rect 1195 29872 1237 29906
rect 1119 29838 1237 29872
rect 1119 29804 1161 29838
rect 1195 29804 1237 29838
rect 1119 29770 1237 29804
rect 1119 29736 1161 29770
rect 1195 29736 1237 29770
rect 1119 29702 1237 29736
rect 1119 29668 1161 29702
rect 1195 29668 1237 29702
rect 1119 29634 1237 29668
rect 1119 29600 1161 29634
rect 1195 29600 1237 29634
rect 1119 29566 1237 29600
rect 1119 29532 1161 29566
rect 1195 29532 1237 29566
rect 1119 29498 1237 29532
rect 1119 29464 1161 29498
rect 1195 29464 1237 29498
rect 1119 29430 1237 29464
rect 1119 29396 1161 29430
rect 1195 29396 1237 29430
rect 1119 29362 1237 29396
rect 1119 29328 1161 29362
rect 1195 29328 1237 29362
rect 1119 29294 1237 29328
rect 1119 29260 1161 29294
rect 1195 29260 1237 29294
rect 1119 29226 1237 29260
rect 1119 29192 1161 29226
rect 1195 29192 1237 29226
rect 1119 29158 1237 29192
rect 1119 29124 1161 29158
rect 1195 29124 1237 29158
rect 1119 29090 1237 29124
rect 1119 29056 1161 29090
rect 1195 29056 1237 29090
rect 1119 29022 1237 29056
rect 1119 28988 1161 29022
rect 1195 28988 1237 29022
rect 1119 28954 1237 28988
rect 1119 28920 1161 28954
rect 1195 28920 1237 28954
rect 1119 28886 1237 28920
rect 13769 34457 13887 34603
rect 13769 34423 13809 34457
rect 13843 34423 13887 34457
rect 13769 34389 13887 34423
rect 13769 34355 13809 34389
rect 13843 34355 13887 34389
rect 13769 34321 13887 34355
rect 13769 34287 13809 34321
rect 13843 34287 13887 34321
rect 13769 34253 13887 34287
rect 13769 34219 13809 34253
rect 13843 34219 13887 34253
rect 13769 34185 13887 34219
rect 13769 34151 13809 34185
rect 13843 34151 13887 34185
rect 13769 34117 13887 34151
rect 13769 34083 13809 34117
rect 13843 34083 13887 34117
rect 13769 34049 13887 34083
rect 13769 34015 13809 34049
rect 13843 34015 13887 34049
rect 13769 33981 13887 34015
rect 13769 33947 13809 33981
rect 13843 33947 13887 33981
rect 13769 33913 13887 33947
rect 13769 33879 13809 33913
rect 13843 33879 13887 33913
rect 13769 33845 13887 33879
rect 13769 33811 13809 33845
rect 13843 33811 13887 33845
rect 13769 33777 13887 33811
rect 13769 33743 13809 33777
rect 13843 33743 13887 33777
rect 13769 33709 13887 33743
rect 13769 33675 13809 33709
rect 13843 33675 13887 33709
rect 13769 33641 13887 33675
rect 13769 33607 13809 33641
rect 13843 33607 13887 33641
rect 13769 33573 13887 33607
rect 13769 33539 13809 33573
rect 13843 33539 13887 33573
rect 13769 33505 13887 33539
rect 13769 33471 13809 33505
rect 13843 33471 13887 33505
rect 13769 33437 13887 33471
rect 13769 33403 13809 33437
rect 13843 33403 13887 33437
rect 13769 33369 13887 33403
rect 13769 33335 13809 33369
rect 13843 33335 13887 33369
rect 13769 33301 13887 33335
rect 13769 33267 13809 33301
rect 13843 33267 13887 33301
rect 13769 33233 13887 33267
rect 13769 33199 13809 33233
rect 13843 33199 13887 33233
rect 13769 33165 13887 33199
rect 13769 33131 13809 33165
rect 13843 33131 13887 33165
rect 13769 33097 13887 33131
rect 13769 33063 13809 33097
rect 13843 33063 13887 33097
rect 13769 33029 13887 33063
rect 13769 32995 13809 33029
rect 13843 32995 13887 33029
rect 13769 32961 13887 32995
rect 13769 32927 13809 32961
rect 13843 32927 13887 32961
rect 13769 32893 13887 32927
rect 13769 32859 13809 32893
rect 13843 32859 13887 32893
rect 13769 32825 13887 32859
rect 13769 32791 13809 32825
rect 13843 32791 13887 32825
rect 13769 32757 13887 32791
rect 13769 32723 13809 32757
rect 13843 32723 13887 32757
rect 13769 32689 13887 32723
rect 13769 32655 13809 32689
rect 13843 32655 13887 32689
rect 13769 32621 13887 32655
rect 13769 32587 13809 32621
rect 13843 32587 13887 32621
rect 13769 32553 13887 32587
rect 13769 32519 13809 32553
rect 13843 32519 13887 32553
rect 13769 32485 13887 32519
rect 13769 32451 13809 32485
rect 13843 32451 13887 32485
rect 13769 32417 13887 32451
rect 13769 32383 13809 32417
rect 13843 32383 13887 32417
rect 13769 32349 13887 32383
rect 13769 32315 13809 32349
rect 13843 32315 13887 32349
rect 13769 32281 13887 32315
rect 13769 32247 13809 32281
rect 13843 32247 13887 32281
rect 13769 32213 13887 32247
rect 13769 32179 13809 32213
rect 13843 32179 13887 32213
rect 13769 32145 13887 32179
rect 13769 32111 13809 32145
rect 13843 32111 13887 32145
rect 13769 32077 13887 32111
rect 13769 32043 13809 32077
rect 13843 32043 13887 32077
rect 13769 32009 13887 32043
rect 13769 31975 13809 32009
rect 13843 31975 13887 32009
rect 13769 31941 13887 31975
rect 13769 31907 13809 31941
rect 13843 31907 13887 31941
rect 13769 31873 13887 31907
rect 13769 31839 13809 31873
rect 13843 31839 13887 31873
rect 13769 31805 13887 31839
rect 13769 31771 13809 31805
rect 13843 31771 13887 31805
rect 13769 31737 13887 31771
rect 13769 31703 13809 31737
rect 13843 31703 13887 31737
rect 13769 31669 13887 31703
rect 13769 31635 13809 31669
rect 13843 31635 13887 31669
rect 13769 31601 13887 31635
rect 13769 31567 13809 31601
rect 13843 31567 13887 31601
rect 13769 31533 13887 31567
rect 13769 31499 13809 31533
rect 13843 31499 13887 31533
rect 13769 31465 13887 31499
rect 13769 31431 13809 31465
rect 13843 31431 13887 31465
rect 13769 31397 13887 31431
rect 13769 31363 13809 31397
rect 13843 31363 13887 31397
rect 13769 31329 13887 31363
rect 13769 31295 13809 31329
rect 13843 31295 13887 31329
rect 13769 31261 13887 31295
rect 13769 31227 13809 31261
rect 13843 31227 13887 31261
rect 13769 31193 13887 31227
rect 13769 31159 13809 31193
rect 13843 31159 13887 31193
rect 13769 31125 13887 31159
rect 13769 31091 13809 31125
rect 13843 31091 13887 31125
rect 13769 31057 13887 31091
rect 13769 31023 13809 31057
rect 13843 31023 13887 31057
rect 13769 30989 13887 31023
rect 13769 30955 13809 30989
rect 13843 30955 13887 30989
rect 13769 30921 13887 30955
rect 13769 30887 13809 30921
rect 13843 30887 13887 30921
rect 13769 30853 13887 30887
rect 13769 30819 13809 30853
rect 13843 30819 13887 30853
rect 13769 30785 13887 30819
rect 13769 30751 13809 30785
rect 13843 30751 13887 30785
rect 13769 30717 13887 30751
rect 13769 30683 13809 30717
rect 13843 30683 13887 30717
rect 13769 30649 13887 30683
rect 13769 30615 13809 30649
rect 13843 30615 13887 30649
rect 13769 30581 13887 30615
rect 13769 30547 13809 30581
rect 13843 30547 13887 30581
rect 13769 30513 13887 30547
rect 13769 30479 13809 30513
rect 13843 30479 13887 30513
rect 13769 30445 13887 30479
rect 13769 30411 13809 30445
rect 13843 30411 13887 30445
rect 13769 30377 13887 30411
rect 13769 30343 13809 30377
rect 13843 30343 13887 30377
rect 13769 30309 13887 30343
rect 13769 30275 13809 30309
rect 13843 30275 13887 30309
rect 13769 30241 13887 30275
rect 13769 30207 13809 30241
rect 13843 30207 13887 30241
rect 13769 30173 13887 30207
rect 13769 30139 13809 30173
rect 13843 30139 13887 30173
rect 13769 30105 13887 30139
rect 13769 30071 13809 30105
rect 13843 30071 13887 30105
rect 13769 30037 13887 30071
rect 13769 30003 13809 30037
rect 13843 30003 13887 30037
rect 13769 29969 13887 30003
rect 13769 29935 13809 29969
rect 13843 29935 13887 29969
rect 13769 29901 13887 29935
rect 13769 29867 13809 29901
rect 13843 29867 13887 29901
rect 13769 29833 13887 29867
rect 13769 29799 13809 29833
rect 13843 29799 13887 29833
rect 13769 29765 13887 29799
rect 13769 29731 13809 29765
rect 13843 29731 13887 29765
rect 13769 29697 13887 29731
rect 13769 29663 13809 29697
rect 13843 29663 13887 29697
rect 13769 29629 13887 29663
rect 13769 29595 13809 29629
rect 13843 29595 13887 29629
rect 13769 29561 13887 29595
rect 13769 29527 13809 29561
rect 13843 29527 13887 29561
rect 13769 29493 13887 29527
rect 13769 29459 13809 29493
rect 13843 29459 13887 29493
rect 13769 29425 13887 29459
rect 13769 29391 13809 29425
rect 13843 29391 13887 29425
rect 13769 29357 13887 29391
rect 13769 29323 13809 29357
rect 13843 29323 13887 29357
rect 13769 29289 13887 29323
rect 13769 29255 13809 29289
rect 13843 29255 13887 29289
rect 13769 29221 13887 29255
rect 13769 29187 13809 29221
rect 13843 29187 13887 29221
rect 13769 29153 13887 29187
rect 13769 29119 13809 29153
rect 13843 29119 13887 29153
rect 13769 29085 13887 29119
rect 13769 29051 13809 29085
rect 13843 29051 13887 29085
rect 13769 29017 13887 29051
rect 13769 28983 13809 29017
rect 13843 28983 13887 29017
rect 13769 28949 13887 28983
rect 13769 28915 13809 28949
rect 13843 28915 13887 28949
rect 1119 28852 1161 28886
rect 1195 28852 1237 28886
rect 1119 28818 1237 28852
rect 1119 28784 1161 28818
rect 1195 28784 1237 28818
rect 1119 28750 1237 28784
rect 1119 28716 1161 28750
rect 1195 28716 1237 28750
rect 1119 28682 1237 28716
rect 1119 28648 1161 28682
rect 1195 28648 1237 28682
rect 1119 28614 1237 28648
rect 1119 28580 1161 28614
rect 1195 28580 1237 28614
rect 1119 28546 1237 28580
rect 1119 28512 1161 28546
rect 1195 28512 1237 28546
rect 1119 28478 1237 28512
rect 1119 28444 1161 28478
rect 1195 28444 1237 28478
rect 1119 28410 1237 28444
rect 1119 28376 1161 28410
rect 1195 28376 1237 28410
rect 1119 28342 1237 28376
rect 1119 28308 1161 28342
rect 1195 28308 1237 28342
rect 1119 28274 1237 28308
rect 1119 28240 1161 28274
rect 1195 28240 1237 28274
rect 1119 28206 1237 28240
rect 1119 28172 1161 28206
rect 1195 28172 1237 28206
rect 1119 28138 1237 28172
rect 1119 28104 1161 28138
rect 1195 28104 1237 28138
rect 1119 28070 1237 28104
rect 1119 28036 1161 28070
rect 1195 28036 1237 28070
rect 1119 28002 1237 28036
rect 1119 27968 1161 28002
rect 1195 27968 1237 28002
rect 1119 27934 1237 27968
rect 1119 27900 1161 27934
rect 1195 27900 1237 27934
rect 1119 27866 1237 27900
rect 1119 27832 1161 27866
rect 1195 27832 1237 27866
rect 1119 27798 1237 27832
rect 1119 27764 1161 27798
rect 1195 27764 1237 27798
rect 1119 27730 1237 27764
rect 1119 27696 1161 27730
rect 1195 27696 1237 27730
rect 1119 27662 1237 27696
rect 1119 27628 1161 27662
rect 1195 27628 1237 27662
rect 1119 27594 1237 27628
rect 1119 27560 1161 27594
rect 1195 27560 1237 27594
rect 1119 27526 1237 27560
rect 1119 27492 1161 27526
rect 1195 27492 1237 27526
rect 1119 27458 1237 27492
rect 1119 27424 1161 27458
rect 1195 27424 1237 27458
rect 1119 27390 1237 27424
rect 1119 27356 1161 27390
rect 1195 27356 1237 27390
rect 1119 27322 1237 27356
rect 1119 27288 1161 27322
rect 1195 27288 1237 27322
rect 1119 27254 1237 27288
rect 1119 27220 1161 27254
rect 1195 27220 1237 27254
rect 1119 27186 1237 27220
rect 1119 27152 1161 27186
rect 1195 27152 1237 27186
rect 1119 27118 1237 27152
rect 1119 27084 1161 27118
rect 1195 27084 1237 27118
rect 1119 27050 1237 27084
rect 1119 27016 1161 27050
rect 1195 27016 1237 27050
rect 13769 28881 13887 28915
rect 13769 28847 13809 28881
rect 13843 28847 13887 28881
rect 13769 28813 13887 28847
rect 13769 28779 13809 28813
rect 13843 28779 13887 28813
rect 13769 28745 13887 28779
rect 13769 28711 13809 28745
rect 13843 28711 13887 28745
rect 13769 28677 13887 28711
rect 13769 28643 13809 28677
rect 13843 28643 13887 28677
rect 13769 28609 13887 28643
rect 13769 28575 13809 28609
rect 13843 28575 13887 28609
rect 13769 28541 13887 28575
rect 13769 28507 13809 28541
rect 13843 28507 13887 28541
rect 13769 28473 13887 28507
rect 13769 28439 13809 28473
rect 13843 28439 13887 28473
rect 13769 28405 13887 28439
rect 13769 28371 13809 28405
rect 13843 28371 13887 28405
rect 13769 28337 13887 28371
rect 13769 28303 13809 28337
rect 13843 28303 13887 28337
rect 13769 28269 13887 28303
rect 13769 28235 13809 28269
rect 13843 28235 13887 28269
rect 13769 28201 13887 28235
rect 13769 28167 13809 28201
rect 13843 28167 13887 28201
rect 13769 28133 13887 28167
rect 13769 28099 13809 28133
rect 13843 28099 13887 28133
rect 13769 28065 13887 28099
rect 13769 28031 13809 28065
rect 13843 28031 13887 28065
rect 13769 27997 13887 28031
rect 13769 27963 13809 27997
rect 13843 27963 13887 27997
rect 13769 27929 13887 27963
rect 13769 27895 13809 27929
rect 13843 27895 13887 27929
rect 13769 27861 13887 27895
rect 13769 27827 13809 27861
rect 13843 27827 13887 27861
rect 13769 27793 13887 27827
rect 13769 27759 13809 27793
rect 13843 27759 13887 27793
rect 13769 27725 13887 27759
rect 13769 27691 13809 27725
rect 13843 27691 13887 27725
rect 13769 27657 13887 27691
rect 13769 27623 13809 27657
rect 13843 27623 13887 27657
rect 13769 27589 13887 27623
rect 13769 27555 13809 27589
rect 13843 27555 13887 27589
rect 13769 27521 13887 27555
rect 13769 27487 13809 27521
rect 13843 27487 13887 27521
rect 13769 27453 13887 27487
rect 13769 27419 13809 27453
rect 13843 27419 13887 27453
rect 13769 27385 13887 27419
rect 13769 27351 13809 27385
rect 13843 27351 13887 27385
rect 13769 27317 13887 27351
rect 13769 27283 13809 27317
rect 13843 27283 13887 27317
rect 13769 27249 13887 27283
rect 13769 27215 13809 27249
rect 13843 27215 13887 27249
rect 13769 27181 13887 27215
rect 13769 27147 13809 27181
rect 13843 27147 13887 27181
rect 13769 27113 13887 27147
rect 13769 27079 13809 27113
rect 13843 27079 13887 27113
rect 13769 27045 13887 27079
rect 1119 26982 1237 27016
rect 1119 26948 1161 26982
rect 1195 26948 1237 26982
rect 1119 26914 1237 26948
rect 1119 26880 1161 26914
rect 1195 26880 1237 26914
rect 1119 26846 1237 26880
rect 1119 26812 1161 26846
rect 1195 26812 1237 26846
rect 1119 26778 1237 26812
rect 1119 26744 1161 26778
rect 1195 26744 1237 26778
rect 1119 26710 1237 26744
rect 1119 26676 1161 26710
rect 1195 26676 1237 26710
rect 1119 26642 1237 26676
rect 1119 26608 1161 26642
rect 1195 26608 1237 26642
rect 1119 26574 1237 26608
rect 1119 26540 1161 26574
rect 1195 26540 1237 26574
rect 1119 26506 1237 26540
rect 1119 26472 1161 26506
rect 1195 26472 1237 26506
rect 1119 26438 1237 26472
rect 1119 26404 1161 26438
rect 1195 26404 1237 26438
rect 1119 26370 1237 26404
rect 1119 26336 1161 26370
rect 1195 26336 1237 26370
rect 1119 26302 1237 26336
rect 1119 26268 1161 26302
rect 1195 26268 1237 26302
rect 1119 26234 1237 26268
rect 1119 26200 1161 26234
rect 1195 26200 1237 26234
rect 1119 26166 1237 26200
rect 1119 26132 1161 26166
rect 1195 26132 1237 26166
rect 1119 26098 1237 26132
rect 1119 26064 1161 26098
rect 1195 26064 1237 26098
rect 1119 26030 1237 26064
rect 1119 25996 1161 26030
rect 1195 25996 1237 26030
rect 1119 25962 1237 25996
rect 1119 25928 1161 25962
rect 1195 25928 1237 25962
rect 1119 25894 1237 25928
rect 1119 25860 1161 25894
rect 1195 25860 1237 25894
rect 1119 25826 1237 25860
rect 1119 25792 1161 25826
rect 1195 25792 1237 25826
rect 1119 25758 1237 25792
rect 1119 25724 1161 25758
rect 1195 25724 1237 25758
rect 1119 25690 1237 25724
rect 1119 25656 1161 25690
rect 1195 25656 1237 25690
rect 1119 25622 1237 25656
rect 1119 25588 1161 25622
rect 1195 25588 1237 25622
rect 1119 25554 1237 25588
rect 1119 25520 1161 25554
rect 1195 25520 1237 25554
rect 1119 25486 1237 25520
rect 1119 25452 1161 25486
rect 1195 25452 1237 25486
rect 1119 25418 1237 25452
rect 1119 25384 1161 25418
rect 1195 25384 1237 25418
rect 1119 25350 1237 25384
rect 1119 25316 1161 25350
rect 1195 25316 1237 25350
rect 1119 25282 1237 25316
rect 1119 25248 1161 25282
rect 1195 25248 1237 25282
rect 1119 25214 1237 25248
rect 1119 25180 1161 25214
rect 1195 25180 1237 25214
rect 1119 25146 1237 25180
rect 1119 25112 1161 25146
rect 1195 25112 1237 25146
rect 1119 25078 1237 25112
rect 1119 25044 1161 25078
rect 1195 25044 1237 25078
rect 1119 25010 1237 25044
rect 1119 24976 1161 25010
rect 1195 24976 1237 25010
rect 1119 24942 1237 24976
rect 1119 24908 1161 24942
rect 1195 24908 1237 24942
rect 1119 24874 1237 24908
rect 1119 24840 1161 24874
rect 1195 24840 1237 24874
rect 1119 24806 1237 24840
rect 1119 24772 1161 24806
rect 1195 24772 1237 24806
rect 1119 24738 1237 24772
rect 1119 24704 1161 24738
rect 1195 24704 1237 24738
rect 1119 24670 1237 24704
rect 1119 24636 1161 24670
rect 1195 24636 1237 24670
rect 1119 24602 1237 24636
rect 1119 24568 1161 24602
rect 1195 24568 1237 24602
rect 1119 24534 1237 24568
rect 1119 24500 1161 24534
rect 1195 24500 1237 24534
rect 1119 24466 1237 24500
rect 1119 24432 1161 24466
rect 1195 24432 1237 24466
rect 1119 24398 1237 24432
rect 1119 24364 1161 24398
rect 1195 24364 1237 24398
rect 1119 24330 1237 24364
rect 1119 24296 1161 24330
rect 1195 24296 1237 24330
rect 1119 24262 1237 24296
rect 1119 24228 1161 24262
rect 1195 24228 1237 24262
rect 1119 24194 1237 24228
rect 1119 24160 1161 24194
rect 1195 24160 1237 24194
rect 1119 24126 1237 24160
rect 1119 24092 1161 24126
rect 1195 24092 1237 24126
rect 1119 24058 1237 24092
rect 1119 24024 1161 24058
rect 1195 24024 1237 24058
rect 1119 23990 1237 24024
rect 1119 23956 1161 23990
rect 1195 23956 1237 23990
rect 1119 23922 1237 23956
rect 1119 23888 1161 23922
rect 1195 23888 1237 23922
rect 1119 23854 1237 23888
rect 1119 23820 1161 23854
rect 1195 23820 1237 23854
rect 1119 23786 1237 23820
rect 1119 23752 1161 23786
rect 1195 23752 1237 23786
rect 1119 23718 1237 23752
rect 1119 23684 1161 23718
rect 1195 23684 1237 23718
rect 1119 23650 1237 23684
rect 1119 23616 1161 23650
rect 1195 23616 1237 23650
rect 1119 23582 1237 23616
rect 1119 23548 1161 23582
rect 1195 23548 1237 23582
rect 1119 23514 1237 23548
rect 1119 23480 1161 23514
rect 1195 23480 1237 23514
rect 1119 23446 1237 23480
rect 1119 23412 1161 23446
rect 1195 23412 1237 23446
rect 1119 23378 1237 23412
rect 1119 23344 1161 23378
rect 1195 23344 1237 23378
rect 1119 23310 1237 23344
rect 1119 23276 1161 23310
rect 1195 23276 1237 23310
rect 1119 23242 1237 23276
rect 1119 23208 1161 23242
rect 1195 23208 1237 23242
rect 1119 23174 1237 23208
rect 1119 23140 1161 23174
rect 1195 23140 1237 23174
rect 1119 23106 1237 23140
rect 1119 23072 1161 23106
rect 1195 23072 1237 23106
rect 1119 23038 1237 23072
rect 1119 23004 1161 23038
rect 1195 23004 1237 23038
rect 1119 22970 1237 23004
rect 1119 22936 1161 22970
rect 1195 22936 1237 22970
rect 1119 22902 1237 22936
rect 1119 22868 1161 22902
rect 1195 22868 1237 22902
rect 1119 22834 1237 22868
rect 1119 22800 1161 22834
rect 1195 22800 1237 22834
rect 1119 22766 1237 22800
rect 1119 22732 1161 22766
rect 1195 22732 1237 22766
rect 1119 22698 1237 22732
rect 1119 22664 1161 22698
rect 1195 22664 1237 22698
rect 1119 22630 1237 22664
rect 1119 22596 1161 22630
rect 1195 22596 1237 22630
rect 1119 22562 1237 22596
rect 1119 22528 1161 22562
rect 1195 22528 1237 22562
rect 1119 22494 1237 22528
rect 1119 22460 1161 22494
rect 1195 22460 1237 22494
rect 1119 22426 1237 22460
rect 1119 22392 1161 22426
rect 1195 22392 1237 22426
rect 1119 22358 1237 22392
rect 1119 22324 1161 22358
rect 1195 22324 1237 22358
rect 1119 22290 1237 22324
rect 1119 22256 1161 22290
rect 1195 22256 1237 22290
rect 1119 22222 1237 22256
rect 1119 22188 1161 22222
rect 1195 22188 1237 22222
rect 1119 22154 1237 22188
rect 1119 22120 1161 22154
rect 1195 22120 1237 22154
rect 1119 22086 1237 22120
rect 1119 22052 1161 22086
rect 1195 22052 1237 22086
rect 1119 22018 1237 22052
rect 1119 21984 1161 22018
rect 1195 21984 1237 22018
rect 1119 21950 1237 21984
rect 1119 21916 1161 21950
rect 1195 21916 1237 21950
rect 1119 21882 1237 21916
rect 1119 21848 1161 21882
rect 1195 21848 1237 21882
rect 1119 21814 1237 21848
rect 1119 21780 1161 21814
rect 1195 21780 1237 21814
rect 1119 21746 1237 21780
rect 1119 21712 1161 21746
rect 1195 21712 1237 21746
rect 1119 21678 1237 21712
rect 1119 21644 1161 21678
rect 1195 21644 1237 21678
rect 1119 21610 1237 21644
rect 1119 21576 1161 21610
rect 1195 21576 1237 21610
rect 1119 21542 1237 21576
rect 1119 21508 1161 21542
rect 1195 21508 1237 21542
rect 1119 21474 1237 21508
rect 1119 21440 1161 21474
rect 1195 21440 1237 21474
rect 1119 21406 1237 21440
rect 1119 21372 1161 21406
rect 1195 21372 1237 21406
rect 1119 21338 1237 21372
rect 1119 21304 1161 21338
rect 1195 21304 1237 21338
rect 1119 21270 1237 21304
rect 1119 21236 1161 21270
rect 1195 21236 1237 21270
rect 1119 21202 1237 21236
rect 1119 21168 1161 21202
rect 1195 21168 1237 21202
rect 1119 21134 1237 21168
rect 1119 21100 1161 21134
rect 1195 21100 1237 21134
rect 1119 21066 1237 21100
rect 1119 21032 1161 21066
rect 1195 21032 1237 21066
rect 1119 20998 1237 21032
rect 1119 20964 1161 20998
rect 1195 20964 1237 20998
rect 1119 20930 1237 20964
rect 1119 20896 1161 20930
rect 1195 20896 1237 20930
rect 1119 20862 1237 20896
rect 1119 20828 1161 20862
rect 1195 20828 1237 20862
rect 1119 20794 1237 20828
rect 1119 20760 1161 20794
rect 1195 20760 1237 20794
rect 1119 20726 1237 20760
rect 1119 20692 1161 20726
rect 1195 20692 1237 20726
rect 1119 20658 1237 20692
rect 1119 20624 1161 20658
rect 1195 20624 1237 20658
rect 1119 20590 1237 20624
rect 1119 20556 1161 20590
rect 1195 20556 1237 20590
rect 1119 20522 1237 20556
rect 1119 20488 1161 20522
rect 1195 20488 1237 20522
rect 1119 20454 1237 20488
rect 1119 20420 1161 20454
rect 1195 20420 1237 20454
rect 1119 20386 1237 20420
rect 1119 20352 1161 20386
rect 1195 20352 1237 20386
rect 1119 20318 1237 20352
rect 1119 20284 1161 20318
rect 1195 20284 1237 20318
rect 1119 20250 1237 20284
rect 1119 20216 1161 20250
rect 1195 20216 1237 20250
rect 1119 20182 1237 20216
rect 1119 20148 1161 20182
rect 1195 20148 1237 20182
rect 1119 20114 1237 20148
rect 1119 20080 1161 20114
rect 1195 20080 1237 20114
rect 1119 20046 1237 20080
rect 1119 20012 1161 20046
rect 1195 20012 1237 20046
rect 1119 19978 1237 20012
rect 1119 19944 1161 19978
rect 1195 19944 1237 19978
rect 1119 19910 1237 19944
rect 1119 19876 1161 19910
rect 1195 19876 1237 19910
rect 1119 19842 1237 19876
rect 1119 19808 1161 19842
rect 1195 19808 1237 19842
rect 1119 19774 1237 19808
rect 1119 19740 1161 19774
rect 1195 19740 1237 19774
rect 1119 19706 1237 19740
rect 1119 19672 1161 19706
rect 1195 19672 1237 19706
rect 1119 19638 1237 19672
rect 1119 19604 1161 19638
rect 1195 19604 1237 19638
rect 1119 19570 1237 19604
rect 1119 19536 1161 19570
rect 1195 19536 1237 19570
rect 1119 19502 1237 19536
rect 1119 19468 1161 19502
rect 1195 19468 1237 19502
rect 1119 19434 1237 19468
rect 1119 19400 1161 19434
rect 1195 19400 1237 19434
rect 1119 19366 1237 19400
rect 1119 19332 1161 19366
rect 1195 19332 1237 19366
rect 1119 19298 1237 19332
rect 1119 19264 1161 19298
rect 1195 19264 1237 19298
rect 1119 19230 1237 19264
rect 1119 19196 1161 19230
rect 1195 19196 1237 19230
rect 1119 19162 1237 19196
rect 1119 19128 1161 19162
rect 1195 19128 1237 19162
rect 1119 19094 1237 19128
rect 1119 19060 1161 19094
rect 1195 19060 1237 19094
rect 1119 19026 1237 19060
rect 1119 18992 1161 19026
rect 1195 18992 1237 19026
rect 1119 18958 1237 18992
rect 1119 18924 1161 18958
rect 1195 18924 1237 18958
rect 1119 18890 1237 18924
rect 1119 18856 1161 18890
rect 1195 18856 1237 18890
rect 1119 18822 1237 18856
rect 1119 18788 1161 18822
rect 1195 18788 1237 18822
rect 1119 18754 1237 18788
rect 1119 18720 1161 18754
rect 1195 18720 1237 18754
rect 1119 18686 1237 18720
rect 1119 18652 1161 18686
rect 1195 18652 1237 18686
rect 1119 18618 1237 18652
rect 1119 18584 1161 18618
rect 1195 18584 1237 18618
rect 1119 18550 1237 18584
rect 1119 18516 1161 18550
rect 1195 18516 1237 18550
rect 1119 18482 1237 18516
rect 1119 18448 1161 18482
rect 1195 18448 1237 18482
rect 1119 18414 1237 18448
rect 1119 18380 1161 18414
rect 1195 18380 1237 18414
rect 1119 18346 1237 18380
rect 1119 18312 1161 18346
rect 1195 18312 1237 18346
rect 1119 18278 1237 18312
rect 1119 18244 1161 18278
rect 1195 18244 1237 18278
rect 1119 18210 1237 18244
rect 1119 18176 1161 18210
rect 1195 18176 1237 18210
rect 1119 18142 1237 18176
rect 1119 18108 1161 18142
rect 1195 18108 1237 18142
rect 1119 18074 1237 18108
rect 1119 18040 1161 18074
rect 1195 18040 1237 18074
rect 1119 18006 1237 18040
rect 1119 17972 1161 18006
rect 1195 17972 1237 18006
rect 1119 17938 1237 17972
rect 1119 17904 1161 17938
rect 1195 17904 1237 17938
rect 1119 17870 1237 17904
rect 1119 17836 1161 17870
rect 1195 17836 1237 17870
rect 1119 17802 1237 17836
rect 1119 17768 1161 17802
rect 1195 17768 1237 17802
rect 1119 17734 1237 17768
rect 1119 17700 1161 17734
rect 1195 17700 1237 17734
rect 1119 17666 1237 17700
rect 1119 17632 1161 17666
rect 1195 17632 1237 17666
rect 1119 17598 1237 17632
rect 1119 17564 1161 17598
rect 1195 17564 1237 17598
rect 1119 17530 1237 17564
rect 1119 17496 1161 17530
rect 1195 17496 1237 17530
rect 1119 17462 1237 17496
rect 1119 17428 1161 17462
rect 1195 17428 1237 17462
rect 1119 17394 1237 17428
rect 1119 17360 1161 17394
rect 1195 17360 1237 17394
rect 1119 17326 1237 17360
rect 1119 17292 1161 17326
rect 1195 17292 1237 17326
rect 1119 17258 1237 17292
rect 1119 17224 1161 17258
rect 1195 17224 1237 17258
rect 1119 17190 1237 17224
rect 1119 17156 1161 17190
rect 1195 17156 1237 17190
rect 1119 17122 1237 17156
rect 1119 17088 1161 17122
rect 1195 17088 1237 17122
rect 1119 17054 1237 17088
rect 1119 17020 1161 17054
rect 1195 17020 1237 17054
rect 1119 16986 1237 17020
rect 1119 16952 1161 16986
rect 1195 16952 1237 16986
rect 1119 16918 1237 16952
rect 1119 16884 1161 16918
rect 1195 16884 1237 16918
rect 1119 16850 1237 16884
rect 1119 16816 1161 16850
rect 1195 16816 1237 16850
rect 1119 16782 1237 16816
rect 1119 16748 1161 16782
rect 1195 16748 1237 16782
rect 1119 16714 1237 16748
rect 1119 16680 1161 16714
rect 1195 16680 1237 16714
rect 1119 16646 1237 16680
rect 1119 16612 1161 16646
rect 1195 16612 1237 16646
rect 1119 16578 1237 16612
rect 1119 16544 1161 16578
rect 1195 16544 1237 16578
rect 1119 16510 1237 16544
rect 1119 16476 1161 16510
rect 1195 16476 1237 16510
rect 1119 16442 1237 16476
rect 1119 16408 1161 16442
rect 1195 16408 1237 16442
rect 1119 16374 1237 16408
rect 1119 16340 1161 16374
rect 1195 16340 1237 16374
rect 1119 16306 1237 16340
rect 1119 16272 1161 16306
rect 1195 16272 1237 16306
rect 1119 16238 1237 16272
rect 1119 16204 1161 16238
rect 1195 16204 1237 16238
rect 1119 16170 1237 16204
rect 1119 16136 1161 16170
rect 1195 16136 1237 16170
rect 1119 16102 1237 16136
rect 1119 16068 1161 16102
rect 1195 16068 1237 16102
rect 1119 16034 1237 16068
rect 1119 16000 1161 16034
rect 1195 16000 1237 16034
rect 1119 15966 1237 16000
rect 1119 15932 1161 15966
rect 1195 15932 1237 15966
rect 1119 15898 1237 15932
rect 1119 15864 1161 15898
rect 1195 15864 1237 15898
rect 1119 15830 1237 15864
rect 1119 15796 1161 15830
rect 1195 15796 1237 15830
rect 1119 15762 1237 15796
rect 1119 15728 1161 15762
rect 1195 15728 1237 15762
rect 1119 15694 1237 15728
rect 1119 15660 1161 15694
rect 1195 15660 1237 15694
rect 1119 15626 1237 15660
rect 1119 15592 1161 15626
rect 1195 15592 1237 15626
rect 1119 15558 1237 15592
rect 1119 15524 1161 15558
rect 1195 15524 1237 15558
rect 1119 15490 1237 15524
rect 1119 15456 1161 15490
rect 1195 15456 1237 15490
rect 1119 15422 1237 15456
rect 1119 15388 1161 15422
rect 1195 15388 1237 15422
rect 1119 15319 1237 15388
rect 13769 27011 13809 27045
rect 13843 27011 13887 27045
rect 13769 26977 13887 27011
rect 13769 26943 13809 26977
rect 13843 26943 13887 26977
rect 13769 26909 13887 26943
rect 13769 26875 13809 26909
rect 13843 26875 13887 26909
rect 13769 26841 13887 26875
rect 13769 26807 13809 26841
rect 13843 26807 13887 26841
rect 13769 26773 13887 26807
rect 13769 26739 13809 26773
rect 13843 26739 13887 26773
rect 13769 26705 13887 26739
rect 13769 26671 13809 26705
rect 13843 26671 13887 26705
rect 13769 26637 13887 26671
rect 13769 26603 13809 26637
rect 13843 26603 13887 26637
rect 13769 26569 13887 26603
rect 13769 26535 13809 26569
rect 13843 26535 13887 26569
rect 13769 26501 13887 26535
rect 13769 26467 13809 26501
rect 13843 26467 13887 26501
rect 13769 26433 13887 26467
rect 13769 26399 13809 26433
rect 13843 26399 13887 26433
rect 13769 26365 13887 26399
rect 13769 26331 13809 26365
rect 13843 26331 13887 26365
rect 13769 26297 13887 26331
rect 13769 26263 13809 26297
rect 13843 26263 13887 26297
rect 13769 26229 13887 26263
rect 13769 26195 13809 26229
rect 13843 26195 13887 26229
rect 13769 26161 13887 26195
rect 13769 26127 13809 26161
rect 13843 26127 13887 26161
rect 13769 26093 13887 26127
rect 13769 26059 13809 26093
rect 13843 26059 13887 26093
rect 13769 26025 13887 26059
rect 13769 25991 13809 26025
rect 13843 25991 13887 26025
rect 13769 25957 13887 25991
rect 13769 25923 13809 25957
rect 13843 25923 13887 25957
rect 13769 25889 13887 25923
rect 13769 25855 13809 25889
rect 13843 25855 13887 25889
rect 13769 25821 13887 25855
rect 13769 25787 13809 25821
rect 13843 25787 13887 25821
rect 13769 25753 13887 25787
rect 13769 25719 13809 25753
rect 13843 25719 13887 25753
rect 13769 25685 13887 25719
rect 13769 25651 13809 25685
rect 13843 25651 13887 25685
rect 13769 25617 13887 25651
rect 13769 25583 13809 25617
rect 13843 25583 13887 25617
rect 13769 25549 13887 25583
rect 13769 25515 13809 25549
rect 13843 25515 13887 25549
rect 13769 25481 13887 25515
rect 13769 25447 13809 25481
rect 13843 25447 13887 25481
rect 13769 25413 13887 25447
rect 13769 25379 13809 25413
rect 13843 25379 13887 25413
rect 13769 25345 13887 25379
rect 13769 25311 13809 25345
rect 13843 25311 13887 25345
rect 13769 25277 13887 25311
rect 13769 25243 13809 25277
rect 13843 25243 13887 25277
rect 13769 25209 13887 25243
rect 13769 25175 13809 25209
rect 13843 25175 13887 25209
rect 13769 25141 13887 25175
rect 13769 25107 13809 25141
rect 13843 25107 13887 25141
rect 13769 25073 13887 25107
rect 13769 25039 13809 25073
rect 13843 25039 13887 25073
rect 13769 25005 13887 25039
rect 13769 24971 13809 25005
rect 13843 24971 13887 25005
rect 13769 24937 13887 24971
rect 13769 24903 13809 24937
rect 13843 24903 13887 24937
rect 13769 24869 13887 24903
rect 13769 24835 13809 24869
rect 13843 24835 13887 24869
rect 13769 24801 13887 24835
rect 13769 24767 13809 24801
rect 13843 24767 13887 24801
rect 13769 24733 13887 24767
rect 13769 24699 13809 24733
rect 13843 24699 13887 24733
rect 13769 24665 13887 24699
rect 13769 24631 13809 24665
rect 13843 24631 13887 24665
rect 13769 24597 13887 24631
rect 13769 24563 13809 24597
rect 13843 24563 13887 24597
rect 13769 24529 13887 24563
rect 13769 24495 13809 24529
rect 13843 24495 13887 24529
rect 13769 24461 13887 24495
rect 13769 24427 13809 24461
rect 13843 24427 13887 24461
rect 13769 24393 13887 24427
rect 13769 24359 13809 24393
rect 13843 24359 13887 24393
rect 13769 24325 13887 24359
rect 13769 24291 13809 24325
rect 13843 24291 13887 24325
rect 13769 24257 13887 24291
rect 13769 24223 13809 24257
rect 13843 24223 13887 24257
rect 13769 24189 13887 24223
rect 13769 24155 13809 24189
rect 13843 24155 13887 24189
rect 13769 24121 13887 24155
rect 13769 24087 13809 24121
rect 13843 24087 13887 24121
rect 13769 24053 13887 24087
rect 13769 24019 13809 24053
rect 13843 24019 13887 24053
rect 13769 23985 13887 24019
rect 13769 23951 13809 23985
rect 13843 23951 13887 23985
rect 13769 23917 13887 23951
rect 13769 23883 13809 23917
rect 13843 23883 13887 23917
rect 13769 23849 13887 23883
rect 13769 23815 13809 23849
rect 13843 23815 13887 23849
rect 13769 23781 13887 23815
rect 13769 23747 13809 23781
rect 13843 23747 13887 23781
rect 13769 23713 13887 23747
rect 13769 23679 13809 23713
rect 13843 23679 13887 23713
rect 13769 23645 13887 23679
rect 13769 23611 13809 23645
rect 13843 23611 13887 23645
rect 13769 23577 13887 23611
rect 13769 23543 13809 23577
rect 13843 23543 13887 23577
rect 13769 23509 13887 23543
rect 13769 23475 13809 23509
rect 13843 23475 13887 23509
rect 13769 23441 13887 23475
rect 13769 23407 13809 23441
rect 13843 23407 13887 23441
rect 13769 23373 13887 23407
rect 13769 23339 13809 23373
rect 13843 23339 13887 23373
rect 13769 23305 13887 23339
rect 13769 23271 13809 23305
rect 13843 23271 13887 23305
rect 13769 23237 13887 23271
rect 13769 23203 13809 23237
rect 13843 23203 13887 23237
rect 13769 23169 13887 23203
rect 13769 23135 13809 23169
rect 13843 23135 13887 23169
rect 13769 23101 13887 23135
rect 13769 23067 13809 23101
rect 13843 23067 13887 23101
rect 13769 23033 13887 23067
rect 13769 22999 13809 23033
rect 13843 22999 13887 23033
rect 13769 22965 13887 22999
rect 13769 22931 13809 22965
rect 13843 22931 13887 22965
rect 13769 22897 13887 22931
rect 13769 22863 13809 22897
rect 13843 22863 13887 22897
rect 13769 22829 13887 22863
rect 13769 22795 13809 22829
rect 13843 22795 13887 22829
rect 13769 22761 13887 22795
rect 13769 22727 13809 22761
rect 13843 22727 13887 22761
rect 13769 22693 13887 22727
rect 13769 22659 13809 22693
rect 13843 22659 13887 22693
rect 13769 22625 13887 22659
rect 13769 22591 13809 22625
rect 13843 22591 13887 22625
rect 13769 22557 13887 22591
rect 13769 22523 13809 22557
rect 13843 22523 13887 22557
rect 13769 22489 13887 22523
rect 13769 22455 13809 22489
rect 13843 22455 13887 22489
rect 13769 22421 13887 22455
rect 13769 22387 13809 22421
rect 13843 22387 13887 22421
rect 13769 22353 13887 22387
rect 13769 22319 13809 22353
rect 13843 22319 13887 22353
rect 13769 22285 13887 22319
rect 13769 22251 13809 22285
rect 13843 22251 13887 22285
rect 13769 22217 13887 22251
rect 13769 22183 13809 22217
rect 13843 22183 13887 22217
rect 13769 22149 13887 22183
rect 13769 22115 13809 22149
rect 13843 22115 13887 22149
rect 13769 22081 13887 22115
rect 13769 22047 13809 22081
rect 13843 22047 13887 22081
rect 13769 22013 13887 22047
rect 13769 21979 13809 22013
rect 13843 21979 13887 22013
rect 13769 21945 13887 21979
rect 13769 21911 13809 21945
rect 13843 21911 13887 21945
rect 13769 21877 13887 21911
rect 13769 21843 13809 21877
rect 13843 21843 13887 21877
rect 13769 21809 13887 21843
rect 13769 21775 13809 21809
rect 13843 21775 13887 21809
rect 13769 21741 13887 21775
rect 13769 21707 13809 21741
rect 13843 21707 13887 21741
rect 13769 21673 13887 21707
rect 13769 21639 13809 21673
rect 13843 21639 13887 21673
rect 13769 21605 13887 21639
rect 13769 21571 13809 21605
rect 13843 21571 13887 21605
rect 13769 21537 13887 21571
rect 13769 21503 13809 21537
rect 13843 21503 13887 21537
rect 13769 21469 13887 21503
rect 13769 21435 13809 21469
rect 13843 21435 13887 21469
rect 13769 21401 13887 21435
rect 13769 21367 13809 21401
rect 13843 21367 13887 21401
rect 13769 21333 13887 21367
rect 13769 21299 13809 21333
rect 13843 21299 13887 21333
rect 13769 21265 13887 21299
rect 13769 21231 13809 21265
rect 13843 21231 13887 21265
rect 13769 21197 13887 21231
rect 13769 21163 13809 21197
rect 13843 21163 13887 21197
rect 13769 21129 13887 21163
rect 13769 21095 13809 21129
rect 13843 21095 13887 21129
rect 13769 21061 13887 21095
rect 13769 21027 13809 21061
rect 13843 21027 13887 21061
rect 13769 20993 13887 21027
rect 13769 20959 13809 20993
rect 13843 20959 13887 20993
rect 13769 20925 13887 20959
rect 13769 20891 13809 20925
rect 13843 20891 13887 20925
rect 13769 20857 13887 20891
rect 13769 20823 13809 20857
rect 13843 20823 13887 20857
rect 13769 20789 13887 20823
rect 13769 20755 13809 20789
rect 13843 20755 13887 20789
rect 13769 20721 13887 20755
rect 13769 20687 13809 20721
rect 13843 20687 13887 20721
rect 13769 20653 13887 20687
rect 13769 20619 13809 20653
rect 13843 20619 13887 20653
rect 13769 20585 13887 20619
rect 13769 20551 13809 20585
rect 13843 20551 13887 20585
rect 13769 20517 13887 20551
rect 13769 20483 13809 20517
rect 13843 20483 13887 20517
rect 13769 20449 13887 20483
rect 13769 20415 13809 20449
rect 13843 20415 13887 20449
rect 13769 20381 13887 20415
rect 13769 20347 13809 20381
rect 13843 20347 13887 20381
rect 13769 20313 13887 20347
rect 13769 20279 13809 20313
rect 13843 20279 13887 20313
rect 13769 20245 13887 20279
rect 13769 20211 13809 20245
rect 13843 20211 13887 20245
rect 13769 20177 13887 20211
rect 13769 20143 13809 20177
rect 13843 20143 13887 20177
rect 13769 20109 13887 20143
rect 13769 20075 13809 20109
rect 13843 20075 13887 20109
rect 13769 20041 13887 20075
rect 13769 20007 13809 20041
rect 13843 20007 13887 20041
rect 13769 19973 13887 20007
rect 13769 19939 13809 19973
rect 13843 19939 13887 19973
rect 13769 19905 13887 19939
rect 13769 19871 13809 19905
rect 13843 19871 13887 19905
rect 13769 19837 13887 19871
rect 13769 19803 13809 19837
rect 13843 19803 13887 19837
rect 13769 19769 13887 19803
rect 13769 19735 13809 19769
rect 13843 19735 13887 19769
rect 13769 19701 13887 19735
rect 13769 19667 13809 19701
rect 13843 19667 13887 19701
rect 13769 19633 13887 19667
rect 13769 19599 13809 19633
rect 13843 19599 13887 19633
rect 13769 19565 13887 19599
rect 13769 19531 13809 19565
rect 13843 19531 13887 19565
rect 13769 19497 13887 19531
rect 13769 19463 13809 19497
rect 13843 19463 13887 19497
rect 13769 19429 13887 19463
rect 13769 19395 13809 19429
rect 13843 19395 13887 19429
rect 13769 19361 13887 19395
rect 13769 19327 13809 19361
rect 13843 19327 13887 19361
rect 13769 19293 13887 19327
rect 13769 19259 13809 19293
rect 13843 19259 13887 19293
rect 13769 19225 13887 19259
rect 13769 19191 13809 19225
rect 13843 19191 13887 19225
rect 13769 19157 13887 19191
rect 13769 19123 13809 19157
rect 13843 19123 13887 19157
rect 13769 19089 13887 19123
rect 13769 19055 13809 19089
rect 13843 19055 13887 19089
rect 13769 19021 13887 19055
rect 13769 18987 13809 19021
rect 13843 18987 13887 19021
rect 13769 18953 13887 18987
rect 13769 18919 13809 18953
rect 13843 18919 13887 18953
rect 13769 18885 13887 18919
rect 13769 18851 13809 18885
rect 13843 18851 13887 18885
rect 13769 18817 13887 18851
rect 13769 18783 13809 18817
rect 13843 18783 13887 18817
rect 13769 18749 13887 18783
rect 13769 18715 13809 18749
rect 13843 18715 13887 18749
rect 13769 18681 13887 18715
rect 13769 18647 13809 18681
rect 13843 18647 13887 18681
rect 13769 18613 13887 18647
rect 13769 18579 13809 18613
rect 13843 18579 13887 18613
rect 13769 18545 13887 18579
rect 13769 18511 13809 18545
rect 13843 18511 13887 18545
rect 13769 18477 13887 18511
rect 13769 18443 13809 18477
rect 13843 18443 13887 18477
rect 13769 18409 13887 18443
rect 13769 18375 13809 18409
rect 13843 18375 13887 18409
rect 13769 18341 13887 18375
rect 13769 18307 13809 18341
rect 13843 18307 13887 18341
rect 13769 18273 13887 18307
rect 13769 18239 13809 18273
rect 13843 18239 13887 18273
rect 13769 18205 13887 18239
rect 13769 18171 13809 18205
rect 13843 18171 13887 18205
rect 13769 18137 13887 18171
rect 13769 18103 13809 18137
rect 13843 18103 13887 18137
rect 13769 18069 13887 18103
rect 13769 18035 13809 18069
rect 13843 18035 13887 18069
rect 13769 18001 13887 18035
rect 13769 17967 13809 18001
rect 13843 17967 13887 18001
rect 13769 17933 13887 17967
rect 13769 17899 13809 17933
rect 13843 17899 13887 17933
rect 13769 17865 13887 17899
rect 13769 17831 13809 17865
rect 13843 17831 13887 17865
rect 13769 17797 13887 17831
rect 13769 17763 13809 17797
rect 13843 17763 13887 17797
rect 13769 17729 13887 17763
rect 13769 17695 13809 17729
rect 13843 17695 13887 17729
rect 13769 17661 13887 17695
rect 13769 17627 13809 17661
rect 13843 17627 13887 17661
rect 13769 17593 13887 17627
rect 13769 17559 13809 17593
rect 13843 17559 13887 17593
rect 13769 17525 13887 17559
rect 13769 17491 13809 17525
rect 13843 17491 13887 17525
rect 13769 17457 13887 17491
rect 13769 17423 13809 17457
rect 13843 17423 13887 17457
rect 13769 17389 13887 17423
rect 13769 17355 13809 17389
rect 13843 17355 13887 17389
rect 13769 17321 13887 17355
rect 13769 17287 13809 17321
rect 13843 17287 13887 17321
rect 13769 17253 13887 17287
rect 13769 17219 13809 17253
rect 13843 17219 13887 17253
rect 13769 17185 13887 17219
rect 13769 17151 13809 17185
rect 13843 17151 13887 17185
rect 13769 17117 13887 17151
rect 13769 17083 13809 17117
rect 13843 17083 13887 17117
rect 13769 17049 13887 17083
rect 13769 17015 13809 17049
rect 13843 17015 13887 17049
rect 13769 16981 13887 17015
rect 13769 16947 13809 16981
rect 13843 16947 13887 16981
rect 13769 16913 13887 16947
rect 13769 16879 13809 16913
rect 13843 16879 13887 16913
rect 13769 16845 13887 16879
rect 13769 16811 13809 16845
rect 13843 16811 13887 16845
rect 13769 16777 13887 16811
rect 13769 16743 13809 16777
rect 13843 16743 13887 16777
rect 13769 16709 13887 16743
rect 13769 16675 13809 16709
rect 13843 16675 13887 16709
rect 13769 16641 13887 16675
rect 13769 16607 13809 16641
rect 13843 16607 13887 16641
rect 13769 16573 13887 16607
rect 13769 16539 13809 16573
rect 13843 16539 13887 16573
rect 13769 16505 13887 16539
rect 13769 16471 13809 16505
rect 13843 16471 13887 16505
rect 13769 16437 13887 16471
rect 13769 16403 13809 16437
rect 13843 16403 13887 16437
rect 13769 16369 13887 16403
rect 13769 16335 13809 16369
rect 13843 16335 13887 16369
rect 13769 16301 13887 16335
rect 13769 16267 13809 16301
rect 13843 16267 13887 16301
rect 13769 16233 13887 16267
rect 13769 16199 13809 16233
rect 13843 16199 13887 16233
rect 13769 16165 13887 16199
rect 13769 16131 13809 16165
rect 13843 16131 13887 16165
rect 13769 16097 13887 16131
rect 13769 16063 13809 16097
rect 13843 16063 13887 16097
rect 13769 16029 13887 16063
rect 13769 15995 13809 16029
rect 13843 15995 13887 16029
rect 13769 15961 13887 15995
rect 13769 15927 13809 15961
rect 13843 15927 13887 15961
rect 13769 15893 13887 15927
rect 13769 15859 13809 15893
rect 13843 15859 13887 15893
rect 13769 15825 13887 15859
rect 13769 15791 13809 15825
rect 13843 15791 13887 15825
rect 13769 15757 13887 15791
rect 13769 15723 13809 15757
rect 13843 15723 13887 15757
rect 13769 15689 13887 15723
rect 13769 15655 13809 15689
rect 13843 15655 13887 15689
rect 13769 15621 13887 15655
rect 13769 15587 13809 15621
rect 13843 15587 13887 15621
rect 13769 15553 13887 15587
rect 13769 15519 13809 15553
rect 13843 15519 13887 15553
rect 13769 15485 13887 15519
rect 13769 15451 13809 15485
rect 13843 15451 13887 15485
rect 13769 15417 13887 15451
rect 13769 15383 13809 15417
rect 13843 15383 13887 15417
rect 13769 15319 13887 15383
rect 1119 15278 13887 15319
rect 1119 15244 1302 15278
rect 1336 15244 1370 15278
rect 1404 15244 1438 15278
rect 1472 15244 1506 15278
rect 1540 15244 1574 15278
rect 1608 15244 1642 15278
rect 1676 15244 1710 15278
rect 1744 15244 1778 15278
rect 1812 15244 1846 15278
rect 1880 15244 1914 15278
rect 1948 15244 1982 15278
rect 2016 15244 2050 15278
rect 2084 15244 2118 15278
rect 2152 15244 2186 15278
rect 2220 15244 2254 15278
rect 2288 15244 2322 15278
rect 2356 15244 2390 15278
rect 2424 15244 2458 15278
rect 2492 15244 2526 15278
rect 2560 15244 2594 15278
rect 2628 15244 2662 15278
rect 2696 15244 2730 15278
rect 2764 15244 2798 15278
rect 2832 15244 2866 15278
rect 2900 15244 2934 15278
rect 2968 15244 3002 15278
rect 3036 15244 3070 15278
rect 3104 15244 3138 15278
rect 3172 15244 3206 15278
rect 3240 15244 3274 15278
rect 3308 15244 3342 15278
rect 3376 15244 3410 15278
rect 3444 15244 3478 15278
rect 3512 15244 3546 15278
rect 3580 15244 3614 15278
rect 3648 15244 3682 15278
rect 3716 15244 3750 15278
rect 3784 15244 3818 15278
rect 3852 15244 3886 15278
rect 3920 15244 3954 15278
rect 3988 15244 4022 15278
rect 4056 15244 4090 15278
rect 4124 15244 4158 15278
rect 4192 15244 4226 15278
rect 4260 15244 4294 15278
rect 4328 15244 4362 15278
rect 4396 15244 4430 15278
rect 4464 15244 4498 15278
rect 4532 15244 4566 15278
rect 4600 15244 4634 15278
rect 4668 15244 4702 15278
rect 4736 15244 4770 15278
rect 4804 15244 4838 15278
rect 4872 15244 4906 15278
rect 4940 15244 4974 15278
rect 5008 15244 5042 15278
rect 5076 15244 5110 15278
rect 5144 15244 5178 15278
rect 5212 15244 5246 15278
rect 5280 15244 5314 15278
rect 5348 15244 5382 15278
rect 5416 15244 5450 15278
rect 5484 15244 5518 15278
rect 5552 15244 5586 15278
rect 5620 15244 5654 15278
rect 5688 15244 5722 15278
rect 5756 15244 5790 15278
rect 5824 15244 5858 15278
rect 5892 15244 5926 15278
rect 5960 15244 5994 15278
rect 6028 15244 6062 15278
rect 6096 15244 6130 15278
rect 6164 15244 6198 15278
rect 6232 15244 6266 15278
rect 6300 15244 6334 15278
rect 6368 15244 6402 15278
rect 6436 15244 6470 15278
rect 6504 15244 6538 15278
rect 6572 15244 6606 15278
rect 6640 15244 6674 15278
rect 6708 15244 6742 15278
rect 6776 15244 6810 15278
rect 6844 15244 6878 15278
rect 6912 15244 6946 15278
rect 6980 15244 7014 15278
rect 7048 15244 7082 15278
rect 7116 15244 7150 15278
rect 7184 15244 7218 15278
rect 7252 15244 7286 15278
rect 7320 15244 7354 15278
rect 7388 15244 7422 15278
rect 7456 15244 7490 15278
rect 7524 15244 7558 15278
rect 7592 15244 7626 15278
rect 7660 15244 7694 15278
rect 7728 15244 7762 15278
rect 7796 15244 7830 15278
rect 7864 15244 7898 15278
rect 7932 15244 7966 15278
rect 8000 15244 8034 15278
rect 8068 15244 8102 15278
rect 8136 15244 8170 15278
rect 8204 15244 8238 15278
rect 8272 15244 8306 15278
rect 8340 15244 8374 15278
rect 8408 15244 8442 15278
rect 8476 15244 8510 15278
rect 8544 15244 8578 15278
rect 8612 15244 8646 15278
rect 8680 15244 8714 15278
rect 8748 15244 8782 15278
rect 8816 15244 8850 15278
rect 8884 15244 8918 15278
rect 8952 15244 8986 15278
rect 9020 15244 9054 15278
rect 9088 15244 9122 15278
rect 9156 15244 9190 15278
rect 9224 15244 9258 15278
rect 9292 15244 9326 15278
rect 9360 15244 9394 15278
rect 9428 15244 9462 15278
rect 9496 15244 9530 15278
rect 9564 15244 9598 15278
rect 9632 15244 9666 15278
rect 9700 15244 9734 15278
rect 9768 15244 9802 15278
rect 9836 15244 9870 15278
rect 9904 15244 9938 15278
rect 9972 15244 10006 15278
rect 10040 15244 10074 15278
rect 10108 15244 10142 15278
rect 10176 15244 10210 15278
rect 10244 15244 10278 15278
rect 10312 15244 10346 15278
rect 10380 15244 10414 15278
rect 10448 15244 10482 15278
rect 10516 15244 10550 15278
rect 10584 15244 10618 15278
rect 10652 15244 10686 15278
rect 10720 15244 10754 15278
rect 10788 15244 10822 15278
rect 10856 15244 10890 15278
rect 10924 15244 10958 15278
rect 10992 15244 11026 15278
rect 11060 15244 11094 15278
rect 11128 15244 11162 15278
rect 11196 15244 11230 15278
rect 11264 15244 11298 15278
rect 11332 15244 11366 15278
rect 11400 15244 11434 15278
rect 11468 15244 11502 15278
rect 11536 15244 11570 15278
rect 11604 15244 11638 15278
rect 11672 15244 11706 15278
rect 11740 15244 11774 15278
rect 11808 15244 11842 15278
rect 11876 15244 11910 15278
rect 11944 15244 11978 15278
rect 12012 15244 12046 15278
rect 12080 15244 12114 15278
rect 12148 15244 12182 15278
rect 12216 15244 12250 15278
rect 12284 15244 12318 15278
rect 12352 15244 12386 15278
rect 12420 15244 12454 15278
rect 12488 15244 12522 15278
rect 12556 15244 12590 15278
rect 12624 15244 12658 15278
rect 12692 15244 12726 15278
rect 12760 15244 12794 15278
rect 12828 15244 12862 15278
rect 12896 15244 12930 15278
rect 12964 15244 12998 15278
rect 13032 15244 13066 15278
rect 13100 15244 13134 15278
rect 13168 15244 13202 15278
rect 13236 15244 13270 15278
rect 13304 15244 13338 15278
rect 13372 15244 13406 15278
rect 13440 15244 13474 15278
rect 13508 15244 13542 15278
rect 13576 15244 13610 15278
rect 13644 15244 13678 15278
rect 13712 15244 13887 15278
rect 1119 15201 13887 15244
rect 14539 36226 14724 36260
rect 14539 36192 14607 36226
rect 14641 36192 14724 36226
rect 14539 36158 14724 36192
rect 14539 36124 14607 36158
rect 14641 36124 14724 36158
rect 14539 36090 14724 36124
rect 14539 36056 14607 36090
rect 14641 36056 14724 36090
rect 14539 36022 14724 36056
rect 14539 35988 14607 36022
rect 14641 35988 14724 36022
rect 14539 35954 14724 35988
rect 14539 35920 14607 35954
rect 14641 35920 14724 35954
rect 14539 35886 14724 35920
rect 14539 35852 14607 35886
rect 14641 35852 14724 35886
rect 14539 35818 14724 35852
rect 14539 35784 14607 35818
rect 14641 35784 14724 35818
rect 14539 35750 14724 35784
rect 14539 35716 14607 35750
rect 14641 35716 14724 35750
rect 14539 35682 14724 35716
rect 14539 35648 14607 35682
rect 14641 35648 14724 35682
rect 14539 35614 14724 35648
rect 14539 35580 14607 35614
rect 14641 35580 14724 35614
rect 14539 35546 14724 35580
rect 14539 35512 14607 35546
rect 14641 35512 14724 35546
rect 14539 35478 14724 35512
rect 14539 35444 14607 35478
rect 14641 35444 14724 35478
rect 14539 35410 14724 35444
rect 14539 35376 14607 35410
rect 14641 35376 14724 35410
rect 14539 35342 14724 35376
rect 14539 35308 14607 35342
rect 14641 35308 14724 35342
rect 14539 35274 14724 35308
rect 14539 35240 14607 35274
rect 14641 35240 14724 35274
rect 14539 35206 14724 35240
rect 14539 35172 14607 35206
rect 14641 35172 14724 35206
rect 14539 35138 14724 35172
rect 14539 35104 14607 35138
rect 14641 35104 14724 35138
rect 14539 35070 14724 35104
rect 14539 35036 14607 35070
rect 14641 35036 14724 35070
rect 14539 35002 14724 35036
rect 14539 34968 14607 35002
rect 14641 34968 14724 35002
rect 14539 34934 14724 34968
rect 14539 34900 14607 34934
rect 14641 34900 14724 34934
rect 14539 34866 14724 34900
rect 14539 34832 14607 34866
rect 14641 34832 14724 34866
rect 14539 34798 14724 34832
rect 14539 34764 14607 34798
rect 14641 34764 14724 34798
rect 14539 34730 14724 34764
rect 14539 34696 14607 34730
rect 14641 34696 14724 34730
rect 14539 34662 14724 34696
rect 14539 34628 14607 34662
rect 14641 34628 14724 34662
rect 14539 34594 14724 34628
rect 14539 34560 14607 34594
rect 14641 34560 14724 34594
rect 14539 34526 14724 34560
rect 14539 34492 14607 34526
rect 14641 34492 14724 34526
rect 14539 34458 14724 34492
rect 14539 34424 14607 34458
rect 14641 34424 14724 34458
rect 14539 34390 14724 34424
rect 14539 34356 14607 34390
rect 14641 34356 14724 34390
rect 14539 34322 14724 34356
rect 14539 34288 14607 34322
rect 14641 34288 14724 34322
rect 14539 34254 14724 34288
rect 14539 34220 14607 34254
rect 14641 34220 14724 34254
rect 14539 34186 14724 34220
rect 14539 34152 14607 34186
rect 14641 34152 14724 34186
rect 14539 34118 14724 34152
rect 14539 34084 14607 34118
rect 14641 34084 14724 34118
rect 14539 34050 14724 34084
rect 14539 34016 14607 34050
rect 14641 34016 14724 34050
rect 14539 33982 14724 34016
rect 14539 33948 14607 33982
rect 14641 33948 14724 33982
rect 14539 33914 14724 33948
rect 14539 33880 14607 33914
rect 14641 33880 14724 33914
rect 14539 33846 14724 33880
rect 14539 33812 14607 33846
rect 14641 33812 14724 33846
rect 14539 33778 14724 33812
rect 14539 33744 14607 33778
rect 14641 33744 14724 33778
rect 14539 33710 14724 33744
rect 14539 33676 14607 33710
rect 14641 33676 14724 33710
rect 14539 33642 14724 33676
rect 14539 33608 14607 33642
rect 14641 33608 14724 33642
rect 14539 33574 14724 33608
rect 14539 33540 14607 33574
rect 14641 33540 14724 33574
rect 14539 33506 14724 33540
rect 14539 33472 14607 33506
rect 14641 33472 14724 33506
rect 14539 33438 14724 33472
rect 14539 33404 14607 33438
rect 14641 33404 14724 33438
rect 14539 33370 14724 33404
rect 14539 33336 14607 33370
rect 14641 33336 14724 33370
rect 14539 33302 14724 33336
rect 14539 33268 14607 33302
rect 14641 33268 14724 33302
rect 14539 33234 14724 33268
rect 14539 33200 14607 33234
rect 14641 33200 14724 33234
rect 14539 33166 14724 33200
rect 14539 33132 14607 33166
rect 14641 33132 14724 33166
rect 14539 33098 14724 33132
rect 14539 33064 14607 33098
rect 14641 33064 14724 33098
rect 14539 33030 14724 33064
rect 14539 32996 14607 33030
rect 14641 32996 14724 33030
rect 14539 32962 14724 32996
rect 14539 32928 14607 32962
rect 14641 32928 14724 32962
rect 14539 32894 14724 32928
rect 14539 32860 14607 32894
rect 14641 32860 14724 32894
rect 14539 32826 14724 32860
rect 14539 32792 14607 32826
rect 14641 32792 14724 32826
rect 14539 32758 14724 32792
rect 14539 32724 14607 32758
rect 14641 32724 14724 32758
rect 14539 32690 14724 32724
rect 14539 32656 14607 32690
rect 14641 32656 14724 32690
rect 14539 32622 14724 32656
rect 14539 32588 14607 32622
rect 14641 32588 14724 32622
rect 14539 32554 14724 32588
rect 14539 32520 14607 32554
rect 14641 32520 14724 32554
rect 14539 32486 14724 32520
rect 14539 32452 14607 32486
rect 14641 32452 14724 32486
rect 14539 32418 14724 32452
rect 14539 32384 14607 32418
rect 14641 32384 14724 32418
rect 14539 32350 14724 32384
rect 14539 32316 14607 32350
rect 14641 32316 14724 32350
rect 14539 32282 14724 32316
rect 14539 32248 14607 32282
rect 14641 32248 14724 32282
rect 14539 32214 14724 32248
rect 14539 32180 14607 32214
rect 14641 32180 14724 32214
rect 14539 32146 14724 32180
rect 14539 32112 14607 32146
rect 14641 32112 14724 32146
rect 14539 32078 14724 32112
rect 14539 32044 14607 32078
rect 14641 32044 14724 32078
rect 14539 32010 14724 32044
rect 14539 31976 14607 32010
rect 14641 31976 14724 32010
rect 14539 31942 14724 31976
rect 14539 31908 14607 31942
rect 14641 31908 14724 31942
rect 14539 31874 14724 31908
rect 14539 31840 14607 31874
rect 14641 31840 14724 31874
rect 14539 31806 14724 31840
rect 14539 31772 14607 31806
rect 14641 31772 14724 31806
rect 14539 31738 14724 31772
rect 14539 31704 14607 31738
rect 14641 31704 14724 31738
rect 14539 31670 14724 31704
rect 14539 31636 14607 31670
rect 14641 31636 14724 31670
rect 14539 31602 14724 31636
rect 14539 31568 14607 31602
rect 14641 31568 14724 31602
rect 14539 31534 14724 31568
rect 14539 31500 14607 31534
rect 14641 31500 14724 31534
rect 14539 31466 14724 31500
rect 14539 31432 14607 31466
rect 14641 31432 14724 31466
rect 14539 31398 14724 31432
rect 14539 31364 14607 31398
rect 14641 31364 14724 31398
rect 14539 31330 14724 31364
rect 14539 31296 14607 31330
rect 14641 31296 14724 31330
rect 14539 31262 14724 31296
rect 14539 31228 14607 31262
rect 14641 31228 14724 31262
rect 14539 31194 14724 31228
rect 14539 31160 14607 31194
rect 14641 31160 14724 31194
rect 14539 31126 14724 31160
rect 14539 31092 14607 31126
rect 14641 31092 14724 31126
rect 14539 31058 14724 31092
rect 14539 31024 14607 31058
rect 14641 31024 14724 31058
rect 14539 30990 14724 31024
rect 14539 30956 14607 30990
rect 14641 30956 14724 30990
rect 14539 30922 14724 30956
rect 14539 30888 14607 30922
rect 14641 30888 14724 30922
rect 14539 30854 14724 30888
rect 14539 30820 14607 30854
rect 14641 30820 14724 30854
rect 14539 30786 14724 30820
rect 14539 30752 14607 30786
rect 14641 30752 14724 30786
rect 14539 30718 14724 30752
rect 14539 30684 14607 30718
rect 14641 30684 14724 30718
rect 14539 30650 14724 30684
rect 14539 30616 14607 30650
rect 14641 30616 14724 30650
rect 14539 30582 14724 30616
rect 14539 30548 14607 30582
rect 14641 30548 14724 30582
rect 14539 30514 14724 30548
rect 14539 30480 14607 30514
rect 14641 30480 14724 30514
rect 14539 30446 14724 30480
rect 14539 30412 14607 30446
rect 14641 30412 14724 30446
rect 14539 30378 14724 30412
rect 14539 30344 14607 30378
rect 14641 30344 14724 30378
rect 14539 30310 14724 30344
rect 14539 30276 14607 30310
rect 14641 30276 14724 30310
rect 14539 30242 14724 30276
rect 14539 30208 14607 30242
rect 14641 30208 14724 30242
rect 14539 30174 14724 30208
rect 14539 30140 14607 30174
rect 14641 30140 14724 30174
rect 14539 30106 14724 30140
rect 14539 30072 14607 30106
rect 14641 30072 14724 30106
rect 14539 30038 14724 30072
rect 14539 30004 14607 30038
rect 14641 30004 14724 30038
rect 14539 29970 14724 30004
rect 14539 29936 14607 29970
rect 14641 29936 14724 29970
rect 14539 29902 14724 29936
rect 14539 29868 14607 29902
rect 14641 29868 14724 29902
rect 14539 29834 14724 29868
rect 14539 29800 14607 29834
rect 14641 29800 14724 29834
rect 14539 29766 14724 29800
rect 14539 29732 14607 29766
rect 14641 29732 14724 29766
rect 14539 29698 14724 29732
rect 14539 29664 14607 29698
rect 14641 29664 14724 29698
rect 14539 29630 14724 29664
rect 14539 29596 14607 29630
rect 14641 29596 14724 29630
rect 14539 29562 14724 29596
rect 14539 29528 14607 29562
rect 14641 29528 14724 29562
rect 14539 29494 14724 29528
rect 14539 29460 14607 29494
rect 14641 29460 14724 29494
rect 14539 29426 14724 29460
rect 14539 29392 14607 29426
rect 14641 29392 14724 29426
rect 14539 29358 14724 29392
rect 14539 29324 14607 29358
rect 14641 29324 14724 29358
rect 14539 29290 14724 29324
rect 14539 29256 14607 29290
rect 14641 29256 14724 29290
rect 14539 29222 14724 29256
rect 14539 29188 14607 29222
rect 14641 29188 14724 29222
rect 14539 29154 14724 29188
rect 14539 29120 14607 29154
rect 14641 29120 14724 29154
rect 14539 29086 14724 29120
rect 14539 29052 14607 29086
rect 14641 29052 14724 29086
rect 14539 29018 14724 29052
rect 14539 28984 14607 29018
rect 14641 28984 14724 29018
rect 14539 28950 14724 28984
rect 14539 28916 14607 28950
rect 14641 28916 14724 28950
rect 14539 28882 14724 28916
rect 14539 28848 14607 28882
rect 14641 28848 14724 28882
rect 14539 28814 14724 28848
rect 14539 28780 14607 28814
rect 14641 28780 14724 28814
rect 14539 28746 14724 28780
rect 14539 28712 14607 28746
rect 14641 28712 14724 28746
rect 14539 28678 14724 28712
rect 14539 28644 14607 28678
rect 14641 28644 14724 28678
rect 14539 28610 14724 28644
rect 14539 28576 14607 28610
rect 14641 28576 14724 28610
rect 14539 28542 14724 28576
rect 14539 28508 14607 28542
rect 14641 28508 14724 28542
rect 14539 28474 14724 28508
rect 14539 28440 14607 28474
rect 14641 28440 14724 28474
rect 14539 28406 14724 28440
rect 14539 28372 14607 28406
rect 14641 28372 14724 28406
rect 14539 28338 14724 28372
rect 14539 28304 14607 28338
rect 14641 28304 14724 28338
rect 14539 28270 14724 28304
rect 14539 28236 14607 28270
rect 14641 28236 14724 28270
rect 14539 28202 14724 28236
rect 14539 28168 14607 28202
rect 14641 28168 14724 28202
rect 14539 28134 14724 28168
rect 14539 28100 14607 28134
rect 14641 28100 14724 28134
rect 14539 28066 14724 28100
rect 14539 28032 14607 28066
rect 14641 28032 14724 28066
rect 14539 27998 14724 28032
rect 14539 27964 14607 27998
rect 14641 27964 14724 27998
rect 14539 27930 14724 27964
rect 14539 27896 14607 27930
rect 14641 27896 14724 27930
rect 14539 27862 14724 27896
rect 14539 27828 14607 27862
rect 14641 27828 14724 27862
rect 14539 27794 14724 27828
rect 14539 27760 14607 27794
rect 14641 27760 14724 27794
rect 14539 27726 14724 27760
rect 14539 27692 14607 27726
rect 14641 27692 14724 27726
rect 14539 27658 14724 27692
rect 14539 27624 14607 27658
rect 14641 27624 14724 27658
rect 14539 27590 14724 27624
rect 14539 27556 14607 27590
rect 14641 27556 14724 27590
rect 14539 27522 14724 27556
rect 14539 27488 14607 27522
rect 14641 27488 14724 27522
rect 14539 27454 14724 27488
rect 14539 27420 14607 27454
rect 14641 27420 14724 27454
rect 14539 27386 14724 27420
rect 14539 27352 14607 27386
rect 14641 27352 14724 27386
rect 14539 27318 14724 27352
rect 14539 27284 14607 27318
rect 14641 27284 14724 27318
rect 14539 27250 14724 27284
rect 14539 27216 14607 27250
rect 14641 27216 14724 27250
rect 14539 27182 14724 27216
rect 14539 27148 14607 27182
rect 14641 27148 14724 27182
rect 14539 27114 14724 27148
rect 14539 27080 14607 27114
rect 14641 27080 14724 27114
rect 14539 27046 14724 27080
rect 14539 27012 14607 27046
rect 14641 27012 14724 27046
rect 14539 26978 14724 27012
rect 14539 26944 14607 26978
rect 14641 26944 14724 26978
rect 14539 26910 14724 26944
rect 14539 26876 14607 26910
rect 14641 26876 14724 26910
rect 14539 26842 14724 26876
rect 14539 26808 14607 26842
rect 14641 26808 14724 26842
rect 14539 26774 14724 26808
rect 14539 26740 14607 26774
rect 14641 26740 14724 26774
rect 14539 26706 14724 26740
rect 14539 26672 14607 26706
rect 14641 26672 14724 26706
rect 14539 26638 14724 26672
rect 14539 26604 14607 26638
rect 14641 26604 14724 26638
rect 14539 26570 14724 26604
rect 14539 26536 14607 26570
rect 14641 26536 14724 26570
rect 14539 26502 14724 26536
rect 14539 26468 14607 26502
rect 14641 26468 14724 26502
rect 14539 26434 14724 26468
rect 14539 26400 14607 26434
rect 14641 26400 14724 26434
rect 14539 26366 14724 26400
rect 14539 26332 14607 26366
rect 14641 26332 14724 26366
rect 14539 26298 14724 26332
rect 14539 26264 14607 26298
rect 14641 26264 14724 26298
rect 14539 26230 14724 26264
rect 14539 26196 14607 26230
rect 14641 26196 14724 26230
rect 14539 26162 14724 26196
rect 14539 26128 14607 26162
rect 14641 26128 14724 26162
rect 14539 26094 14724 26128
rect 14539 26060 14607 26094
rect 14641 26060 14724 26094
rect 14539 26026 14724 26060
rect 14539 25992 14607 26026
rect 14641 25992 14724 26026
rect 14539 25958 14724 25992
rect 14539 25924 14607 25958
rect 14641 25924 14724 25958
rect 14539 25890 14724 25924
rect 14539 25856 14607 25890
rect 14641 25856 14724 25890
rect 14539 25822 14724 25856
rect 14539 25788 14607 25822
rect 14641 25788 14724 25822
rect 14539 25754 14724 25788
rect 14539 25720 14607 25754
rect 14641 25720 14724 25754
rect 14539 25686 14724 25720
rect 14539 25652 14607 25686
rect 14641 25652 14724 25686
rect 14539 25618 14724 25652
rect 14539 25584 14607 25618
rect 14641 25584 14724 25618
rect 14539 25550 14724 25584
rect 14539 25516 14607 25550
rect 14641 25516 14724 25550
rect 14539 25482 14724 25516
rect 14539 25448 14607 25482
rect 14641 25448 14724 25482
rect 14539 25414 14724 25448
rect 14539 25380 14607 25414
rect 14641 25380 14724 25414
rect 14539 25346 14724 25380
rect 14539 25312 14607 25346
rect 14641 25312 14724 25346
rect 14539 25278 14724 25312
rect 14539 25244 14607 25278
rect 14641 25244 14724 25278
rect 14539 25210 14724 25244
rect 14539 25176 14607 25210
rect 14641 25176 14724 25210
rect 14539 25142 14724 25176
rect 14539 25108 14607 25142
rect 14641 25108 14724 25142
rect 14539 25074 14724 25108
rect 14539 25040 14607 25074
rect 14641 25040 14724 25074
rect 14539 25006 14724 25040
rect 14539 24972 14607 25006
rect 14641 24972 14724 25006
rect 14539 24938 14724 24972
rect 14539 24904 14607 24938
rect 14641 24904 14724 24938
rect 14539 24870 14724 24904
rect 14539 24836 14607 24870
rect 14641 24836 14724 24870
rect 14539 24802 14724 24836
rect 14539 24768 14607 24802
rect 14641 24768 14724 24802
rect 14539 24734 14724 24768
rect 14539 24700 14607 24734
rect 14641 24700 14724 24734
rect 14539 24666 14724 24700
rect 14539 24632 14607 24666
rect 14641 24632 14724 24666
rect 14539 24598 14724 24632
rect 14539 24564 14607 24598
rect 14641 24564 14724 24598
rect 14539 24530 14724 24564
rect 14539 24496 14607 24530
rect 14641 24496 14724 24530
rect 14539 24462 14724 24496
rect 14539 24428 14607 24462
rect 14641 24428 14724 24462
rect 14539 24394 14724 24428
rect 14539 24360 14607 24394
rect 14641 24360 14724 24394
rect 14539 24326 14724 24360
rect 14539 24292 14607 24326
rect 14641 24292 14724 24326
rect 14539 24258 14724 24292
rect 14539 24224 14607 24258
rect 14641 24224 14724 24258
rect 14539 24190 14724 24224
rect 14539 24156 14607 24190
rect 14641 24156 14724 24190
rect 14539 24122 14724 24156
rect 14539 24088 14607 24122
rect 14641 24088 14724 24122
rect 14539 24054 14724 24088
rect 14539 24020 14607 24054
rect 14641 24020 14724 24054
rect 14539 23986 14724 24020
rect 14539 23952 14607 23986
rect 14641 23952 14724 23986
rect 14539 23918 14724 23952
rect 14539 23884 14607 23918
rect 14641 23884 14724 23918
rect 14539 23850 14724 23884
rect 14539 23816 14607 23850
rect 14641 23816 14724 23850
rect 14539 23782 14724 23816
rect 14539 23748 14607 23782
rect 14641 23748 14724 23782
rect 14539 23714 14724 23748
rect 14539 23680 14607 23714
rect 14641 23680 14724 23714
rect 14539 23646 14724 23680
rect 14539 23612 14607 23646
rect 14641 23612 14724 23646
rect 14539 23578 14724 23612
rect 14539 23544 14607 23578
rect 14641 23544 14724 23578
rect 14539 23510 14724 23544
rect 14539 23476 14607 23510
rect 14641 23476 14724 23510
rect 14539 23442 14724 23476
rect 14539 23408 14607 23442
rect 14641 23408 14724 23442
rect 14539 23374 14724 23408
rect 14539 23340 14607 23374
rect 14641 23340 14724 23374
rect 14539 23306 14724 23340
rect 14539 23272 14607 23306
rect 14641 23272 14724 23306
rect 14539 23238 14724 23272
rect 14539 23204 14607 23238
rect 14641 23204 14724 23238
rect 14539 23170 14724 23204
rect 14539 23136 14607 23170
rect 14641 23136 14724 23170
rect 14539 23102 14724 23136
rect 14539 23068 14607 23102
rect 14641 23068 14724 23102
rect 14539 23034 14724 23068
rect 14539 23000 14607 23034
rect 14641 23000 14724 23034
rect 14539 22966 14724 23000
rect 14539 22932 14607 22966
rect 14641 22932 14724 22966
rect 14539 22898 14724 22932
rect 14539 22864 14607 22898
rect 14641 22864 14724 22898
rect 14539 22830 14724 22864
rect 14539 22796 14607 22830
rect 14641 22796 14724 22830
rect 14539 22762 14724 22796
rect 14539 22728 14607 22762
rect 14641 22728 14724 22762
rect 14539 22694 14724 22728
rect 14539 22660 14607 22694
rect 14641 22660 14724 22694
rect 14539 22626 14724 22660
rect 14539 22592 14607 22626
rect 14641 22592 14724 22626
rect 14539 22558 14724 22592
rect 14539 22524 14607 22558
rect 14641 22524 14724 22558
rect 14539 22490 14724 22524
rect 14539 22456 14607 22490
rect 14641 22456 14724 22490
rect 14539 22422 14724 22456
rect 14539 22388 14607 22422
rect 14641 22388 14724 22422
rect 14539 22354 14724 22388
rect 14539 22320 14607 22354
rect 14641 22320 14724 22354
rect 14539 22286 14724 22320
rect 14539 22252 14607 22286
rect 14641 22252 14724 22286
rect 14539 22218 14724 22252
rect 14539 22184 14607 22218
rect 14641 22184 14724 22218
rect 14539 22150 14724 22184
rect 14539 22116 14607 22150
rect 14641 22116 14724 22150
rect 14539 22082 14724 22116
rect 14539 22048 14607 22082
rect 14641 22048 14724 22082
rect 14539 22014 14724 22048
rect 14539 21980 14607 22014
rect 14641 21980 14724 22014
rect 14539 21946 14724 21980
rect 14539 21912 14607 21946
rect 14641 21912 14724 21946
rect 14539 21878 14724 21912
rect 14539 21844 14607 21878
rect 14641 21844 14724 21878
rect 14539 21810 14724 21844
rect 14539 21776 14607 21810
rect 14641 21776 14724 21810
rect 14539 21742 14724 21776
rect 14539 21708 14607 21742
rect 14641 21708 14724 21742
rect 14539 21674 14724 21708
rect 14539 21640 14607 21674
rect 14641 21640 14724 21674
rect 14539 21606 14724 21640
rect 14539 21572 14607 21606
rect 14641 21572 14724 21606
rect 14539 21538 14724 21572
rect 14539 21504 14607 21538
rect 14641 21504 14724 21538
rect 14539 21470 14724 21504
rect 14539 21436 14607 21470
rect 14641 21436 14724 21470
rect 14539 21402 14724 21436
rect 14539 21368 14607 21402
rect 14641 21368 14724 21402
rect 14539 21334 14724 21368
rect 14539 21300 14607 21334
rect 14641 21300 14724 21334
rect 14539 21266 14724 21300
rect 14539 21232 14607 21266
rect 14641 21232 14724 21266
rect 14539 21198 14724 21232
rect 14539 21164 14607 21198
rect 14641 21164 14724 21198
rect 14539 21130 14724 21164
rect 14539 21096 14607 21130
rect 14641 21096 14724 21130
rect 14539 21062 14724 21096
rect 14539 21028 14607 21062
rect 14641 21028 14724 21062
rect 14539 20994 14724 21028
rect 14539 20960 14607 20994
rect 14641 20960 14724 20994
rect 14539 20926 14724 20960
rect 14539 20892 14607 20926
rect 14641 20892 14724 20926
rect 14539 20858 14724 20892
rect 14539 20824 14607 20858
rect 14641 20824 14724 20858
rect 14539 20790 14724 20824
rect 14539 20756 14607 20790
rect 14641 20756 14724 20790
rect 14539 20722 14724 20756
rect 14539 20688 14607 20722
rect 14641 20688 14724 20722
rect 14539 20654 14724 20688
rect 14539 20620 14607 20654
rect 14641 20620 14724 20654
rect 14539 20586 14724 20620
rect 14539 20552 14607 20586
rect 14641 20552 14724 20586
rect 14539 20518 14724 20552
rect 14539 20484 14607 20518
rect 14641 20484 14724 20518
rect 14539 20450 14724 20484
rect 14539 20416 14607 20450
rect 14641 20416 14724 20450
rect 14539 20382 14724 20416
rect 14539 20348 14607 20382
rect 14641 20348 14724 20382
rect 14539 20314 14724 20348
rect 14539 20280 14607 20314
rect 14641 20280 14724 20314
rect 14539 20246 14724 20280
rect 14539 20212 14607 20246
rect 14641 20212 14724 20246
rect 14539 20178 14724 20212
rect 14539 20144 14607 20178
rect 14641 20144 14724 20178
rect 14539 20110 14724 20144
rect 14539 20076 14607 20110
rect 14641 20076 14724 20110
rect 14539 20042 14724 20076
rect 14539 20008 14607 20042
rect 14641 20008 14724 20042
rect 14539 19974 14724 20008
rect 14539 19940 14607 19974
rect 14641 19940 14724 19974
rect 14539 19906 14724 19940
rect 14539 19872 14607 19906
rect 14641 19872 14724 19906
rect 14539 19838 14724 19872
rect 14539 19804 14607 19838
rect 14641 19804 14724 19838
rect 14539 19770 14724 19804
rect 14539 19736 14607 19770
rect 14641 19736 14724 19770
rect 14539 19702 14724 19736
rect 14539 19668 14607 19702
rect 14641 19668 14724 19702
rect 14539 19634 14724 19668
rect 14539 19600 14607 19634
rect 14641 19600 14724 19634
rect 14539 19566 14724 19600
rect 14539 19532 14607 19566
rect 14641 19532 14724 19566
rect 14539 19498 14724 19532
rect 14539 19464 14607 19498
rect 14641 19464 14724 19498
rect 14539 19430 14724 19464
rect 14539 19396 14607 19430
rect 14641 19396 14724 19430
rect 14539 19362 14724 19396
rect 14539 19328 14607 19362
rect 14641 19328 14724 19362
rect 14539 19294 14724 19328
rect 14539 19260 14607 19294
rect 14641 19260 14724 19294
rect 14539 19226 14724 19260
rect 14539 19192 14607 19226
rect 14641 19192 14724 19226
rect 14539 19158 14724 19192
rect 14539 19124 14607 19158
rect 14641 19124 14724 19158
rect 14539 19090 14724 19124
rect 14539 19056 14607 19090
rect 14641 19056 14724 19090
rect 14539 19022 14724 19056
rect 14539 18988 14607 19022
rect 14641 18988 14724 19022
rect 14539 18954 14724 18988
rect 14539 18920 14607 18954
rect 14641 18920 14724 18954
rect 14539 18886 14724 18920
rect 14539 18852 14607 18886
rect 14641 18852 14724 18886
rect 14539 18818 14724 18852
rect 14539 18784 14607 18818
rect 14641 18784 14724 18818
rect 14539 18750 14724 18784
rect 14539 18716 14607 18750
rect 14641 18716 14724 18750
rect 14539 18682 14724 18716
rect 14539 18648 14607 18682
rect 14641 18648 14724 18682
rect 14539 18614 14724 18648
rect 14539 18580 14607 18614
rect 14641 18580 14724 18614
rect 14539 18546 14724 18580
rect 14539 18512 14607 18546
rect 14641 18512 14724 18546
rect 14539 18478 14724 18512
rect 14539 18444 14607 18478
rect 14641 18444 14724 18478
rect 14539 18410 14724 18444
rect 14539 18376 14607 18410
rect 14641 18376 14724 18410
rect 14539 18342 14724 18376
rect 14539 18308 14607 18342
rect 14641 18308 14724 18342
rect 14539 18274 14724 18308
rect 14539 18240 14607 18274
rect 14641 18240 14724 18274
rect 14539 18206 14724 18240
rect 14539 18172 14607 18206
rect 14641 18172 14724 18206
rect 14539 18138 14724 18172
rect 14539 18104 14607 18138
rect 14641 18104 14724 18138
rect 14539 18070 14724 18104
rect 14539 18036 14607 18070
rect 14641 18036 14724 18070
rect 14539 18002 14724 18036
rect 14539 17968 14607 18002
rect 14641 17968 14724 18002
rect 14539 17934 14724 17968
rect 14539 17900 14607 17934
rect 14641 17900 14724 17934
rect 14539 17866 14724 17900
rect 14539 17832 14607 17866
rect 14641 17832 14724 17866
rect 14539 17798 14724 17832
rect 14539 17764 14607 17798
rect 14641 17764 14724 17798
rect 14539 17730 14724 17764
rect 14539 17696 14607 17730
rect 14641 17696 14724 17730
rect 14539 17662 14724 17696
rect 14539 17628 14607 17662
rect 14641 17628 14724 17662
rect 14539 17594 14724 17628
rect 14539 17560 14607 17594
rect 14641 17560 14724 17594
rect 14539 17526 14724 17560
rect 14539 17492 14607 17526
rect 14641 17492 14724 17526
rect 14539 17458 14724 17492
rect 14539 17424 14607 17458
rect 14641 17424 14724 17458
rect 14539 17390 14724 17424
rect 14539 17356 14607 17390
rect 14641 17356 14724 17390
rect 14539 17322 14724 17356
rect 14539 17288 14607 17322
rect 14641 17288 14724 17322
rect 14539 17254 14724 17288
rect 14539 17220 14607 17254
rect 14641 17220 14724 17254
rect 14539 17186 14724 17220
rect 14539 17152 14607 17186
rect 14641 17152 14724 17186
rect 14539 17118 14724 17152
rect 14539 17084 14607 17118
rect 14641 17084 14724 17118
rect 14539 17050 14724 17084
rect 14539 17016 14607 17050
rect 14641 17016 14724 17050
rect 14539 16982 14724 17016
rect 14539 16948 14607 16982
rect 14641 16948 14724 16982
rect 14539 16914 14724 16948
rect 14539 16880 14607 16914
rect 14641 16880 14724 16914
rect 14539 16846 14724 16880
rect 14539 16812 14607 16846
rect 14641 16812 14724 16846
rect 14539 16778 14724 16812
rect 14539 16744 14607 16778
rect 14641 16744 14724 16778
rect 14539 16710 14724 16744
rect 14539 16676 14607 16710
rect 14641 16676 14724 16710
rect 14539 16642 14724 16676
rect 14539 16608 14607 16642
rect 14641 16608 14724 16642
rect 14539 16574 14724 16608
rect 14539 16540 14607 16574
rect 14641 16540 14724 16574
rect 14539 16506 14724 16540
rect 14539 16472 14607 16506
rect 14641 16472 14724 16506
rect 14539 16438 14724 16472
rect 14539 16404 14607 16438
rect 14641 16404 14724 16438
rect 14539 16370 14724 16404
rect 14539 16336 14607 16370
rect 14641 16336 14724 16370
rect 14539 16302 14724 16336
rect 14539 16268 14607 16302
rect 14641 16268 14724 16302
rect 14539 16234 14724 16268
rect 14539 16200 14607 16234
rect 14641 16200 14724 16234
rect 14539 16166 14724 16200
rect 14539 16132 14607 16166
rect 14641 16132 14724 16166
rect 14539 16098 14724 16132
rect 14539 16064 14607 16098
rect 14641 16064 14724 16098
rect 14539 16030 14724 16064
rect 14539 15996 14607 16030
rect 14641 15996 14724 16030
rect 14539 15962 14724 15996
rect 14539 15928 14607 15962
rect 14641 15928 14724 15962
rect 14539 15894 14724 15928
rect 14539 15860 14607 15894
rect 14641 15860 14724 15894
rect 14539 15826 14724 15860
rect 14539 15792 14607 15826
rect 14641 15792 14724 15826
rect 14539 15758 14724 15792
rect 14539 15724 14607 15758
rect 14641 15724 14724 15758
rect 14539 15690 14724 15724
rect 14539 15656 14607 15690
rect 14641 15656 14724 15690
rect 14539 15622 14724 15656
rect 14539 15588 14607 15622
rect 14641 15588 14724 15622
rect 14539 15554 14724 15588
rect 14539 15520 14607 15554
rect 14641 15520 14724 15554
rect 14539 15486 14724 15520
rect 14539 15452 14607 15486
rect 14641 15452 14724 15486
rect 14539 15418 14724 15452
rect 14539 15384 14607 15418
rect 14641 15384 14724 15418
rect 14539 15350 14724 15384
rect 14539 15316 14607 15350
rect 14641 15316 14724 15350
rect 14539 15282 14724 15316
rect 14539 15248 14607 15282
rect 14641 15248 14724 15282
rect 14539 15214 14724 15248
rect 14539 15180 14607 15214
rect 14641 15180 14724 15214
rect 14539 15146 14724 15180
rect 14539 15112 14607 15146
rect 14641 15112 14724 15146
rect 14539 15078 14724 15112
rect 14539 15044 14607 15078
rect 14641 15044 14724 15078
rect 14539 15010 14724 15044
rect 14539 14976 14607 15010
rect 14641 14976 14724 15010
rect 14539 14942 14724 14976
rect 14539 14908 14607 14942
rect 14641 14908 14724 14942
rect 14539 14874 14724 14908
rect 14539 14840 14607 14874
rect 14641 14840 14724 14874
rect 14539 14806 14724 14840
rect 14539 14772 14607 14806
rect 14641 14772 14724 14806
rect 14539 14738 14724 14772
rect 14539 14704 14607 14738
rect 14641 14704 14724 14738
rect 245 14630 312 14664
rect 346 14630 430 14664
rect 245 14596 430 14630
rect 245 14562 312 14596
rect 346 14562 430 14596
rect 245 14528 430 14562
rect 14539 14670 14724 14704
rect 14539 14636 14607 14670
rect 14641 14636 14724 14670
rect 14539 14602 14724 14636
rect 14539 14568 14607 14602
rect 14641 14568 14724 14602
rect 14539 14528 14724 14568
rect 245 14451 14724 14528
rect 245 14417 476 14451
rect 510 14417 544 14451
rect 578 14417 612 14451
rect 646 14417 680 14451
rect 714 14417 748 14451
rect 782 14417 816 14451
rect 850 14417 884 14451
rect 918 14417 952 14451
rect 986 14417 1020 14451
rect 1054 14417 1088 14451
rect 1122 14417 1156 14451
rect 1190 14417 1224 14451
rect 1258 14417 1292 14451
rect 1326 14417 1360 14451
rect 1394 14417 1428 14451
rect 1462 14417 1496 14451
rect 1530 14417 1564 14451
rect 1598 14417 1632 14451
rect 1666 14417 1700 14451
rect 1734 14417 1768 14451
rect 1802 14417 1836 14451
rect 1870 14417 1904 14451
rect 1938 14417 1972 14451
rect 2006 14417 2040 14451
rect 2074 14417 2108 14451
rect 2142 14417 2176 14451
rect 2210 14417 2244 14451
rect 2278 14417 2312 14451
rect 2346 14417 2380 14451
rect 2414 14417 2448 14451
rect 2482 14417 2516 14451
rect 2550 14417 2584 14451
rect 2618 14417 2652 14451
rect 2686 14417 2720 14451
rect 2754 14417 2788 14451
rect 2822 14417 2856 14451
rect 2890 14417 2924 14451
rect 2958 14417 2992 14451
rect 3026 14417 3060 14451
rect 3094 14417 3128 14451
rect 3162 14417 3196 14451
rect 3230 14417 3264 14451
rect 3298 14417 3332 14451
rect 3366 14417 3400 14451
rect 3434 14417 3468 14451
rect 3502 14417 3536 14451
rect 3570 14417 3604 14451
rect 3638 14417 3672 14451
rect 3706 14417 3740 14451
rect 3774 14417 3808 14451
rect 3842 14417 3876 14451
rect 3910 14417 3944 14451
rect 3978 14417 4012 14451
rect 4046 14417 4080 14451
rect 4114 14417 4148 14451
rect 4182 14417 4216 14451
rect 4250 14417 4284 14451
rect 4318 14417 4352 14451
rect 4386 14417 4420 14451
rect 4454 14417 4488 14451
rect 4522 14417 4556 14451
rect 4590 14417 4624 14451
rect 4658 14417 4692 14451
rect 4726 14417 4760 14451
rect 4794 14417 4828 14451
rect 4862 14417 4896 14451
rect 4930 14417 4964 14451
rect 4998 14417 5032 14451
rect 5066 14417 5100 14451
rect 5134 14417 5168 14451
rect 5202 14417 5236 14451
rect 5270 14417 5304 14451
rect 5338 14417 5372 14451
rect 5406 14417 5440 14451
rect 5474 14417 5508 14451
rect 5542 14417 5576 14451
rect 5610 14417 5644 14451
rect 5678 14417 5712 14451
rect 5746 14417 5780 14451
rect 5814 14417 5848 14451
rect 5882 14417 5916 14451
rect 5950 14417 5984 14451
rect 6018 14417 6052 14451
rect 6086 14417 6120 14451
rect 6154 14417 6188 14451
rect 6222 14417 6256 14451
rect 6290 14417 6324 14451
rect 6358 14417 6392 14451
rect 6426 14417 6460 14451
rect 6494 14417 6528 14451
rect 6562 14417 6596 14451
rect 6630 14417 6664 14451
rect 6698 14417 6732 14451
rect 6766 14417 6800 14451
rect 6834 14417 6868 14451
rect 6902 14417 6936 14451
rect 6970 14417 7004 14451
rect 7038 14417 7072 14451
rect 7106 14417 7140 14451
rect 7174 14417 7208 14451
rect 7242 14417 7276 14451
rect 7310 14417 7344 14451
rect 7378 14417 7412 14451
rect 7446 14417 7480 14451
rect 7514 14417 7548 14451
rect 7582 14417 7616 14451
rect 7650 14417 7684 14451
rect 7718 14417 7752 14451
rect 7786 14417 7820 14451
rect 7854 14417 7888 14451
rect 7922 14417 7956 14451
rect 7990 14417 8024 14451
rect 8058 14417 8092 14451
rect 8126 14417 8160 14451
rect 8194 14417 8228 14451
rect 8262 14417 8296 14451
rect 8330 14417 8364 14451
rect 8398 14417 8432 14451
rect 8466 14417 8500 14451
rect 8534 14417 8568 14451
rect 8602 14417 8636 14451
rect 8670 14417 8704 14451
rect 8738 14417 8772 14451
rect 8806 14417 8840 14451
rect 8874 14417 8908 14451
rect 8942 14417 8976 14451
rect 9010 14417 9044 14451
rect 9078 14417 9112 14451
rect 9146 14417 9180 14451
rect 9214 14417 9248 14451
rect 9282 14417 9316 14451
rect 9350 14417 9384 14451
rect 9418 14417 9452 14451
rect 9486 14417 9520 14451
rect 9554 14417 9588 14451
rect 9622 14417 9656 14451
rect 9690 14417 9724 14451
rect 9758 14417 9792 14451
rect 9826 14417 9860 14451
rect 9894 14417 9928 14451
rect 9962 14417 9996 14451
rect 10030 14417 10064 14451
rect 10098 14417 10132 14451
rect 10166 14417 10200 14451
rect 10234 14417 10268 14451
rect 10302 14417 10336 14451
rect 10370 14417 10404 14451
rect 10438 14417 10472 14451
rect 10506 14417 10540 14451
rect 10574 14417 10608 14451
rect 10642 14417 10676 14451
rect 10710 14417 10744 14451
rect 10778 14417 10812 14451
rect 10846 14417 10880 14451
rect 10914 14417 10948 14451
rect 10982 14417 11016 14451
rect 11050 14417 11084 14451
rect 11118 14417 11152 14451
rect 11186 14417 11220 14451
rect 11254 14417 11288 14451
rect 11322 14417 11356 14451
rect 11390 14417 11424 14451
rect 11458 14417 11492 14451
rect 11526 14417 11560 14451
rect 11594 14417 11628 14451
rect 11662 14417 11696 14451
rect 11730 14417 11764 14451
rect 11798 14417 11832 14451
rect 11866 14417 11900 14451
rect 11934 14417 11968 14451
rect 12002 14417 12036 14451
rect 12070 14417 12104 14451
rect 12138 14417 12172 14451
rect 12206 14417 12240 14451
rect 12274 14417 12308 14451
rect 12342 14417 12376 14451
rect 12410 14417 12444 14451
rect 12478 14417 12512 14451
rect 12546 14417 12580 14451
rect 12614 14417 12648 14451
rect 12682 14417 12716 14451
rect 12750 14417 12784 14451
rect 12818 14417 12852 14451
rect 12886 14417 12920 14451
rect 12954 14417 12988 14451
rect 13022 14417 13056 14451
rect 13090 14417 13124 14451
rect 13158 14417 13192 14451
rect 13226 14417 13260 14451
rect 13294 14417 13328 14451
rect 13362 14417 13396 14451
rect 13430 14417 13464 14451
rect 13498 14417 13532 14451
rect 13566 14417 13600 14451
rect 13634 14417 13668 14451
rect 13702 14417 13736 14451
rect 13770 14417 13804 14451
rect 13838 14417 13872 14451
rect 13906 14417 13940 14451
rect 13974 14417 14008 14451
rect 14042 14417 14076 14451
rect 14110 14417 14144 14451
rect 14178 14417 14212 14451
rect 14246 14417 14280 14451
rect 14314 14417 14348 14451
rect 14382 14417 14416 14451
rect 14450 14417 14484 14451
rect 14518 14417 14724 14451
rect 245 14343 14724 14417
<< mvnsubdiff >>
rect 583 36177 14381 36227
rect 583 36143 766 36177
rect 800 36143 834 36177
rect 868 36143 902 36177
rect 936 36143 970 36177
rect 1004 36143 1038 36177
rect 1072 36143 1106 36177
rect 1140 36143 1174 36177
rect 1208 36143 1242 36177
rect 1276 36143 1310 36177
rect 1344 36143 1378 36177
rect 1412 36143 1446 36177
rect 1480 36143 1514 36177
rect 1548 36143 1582 36177
rect 1616 36143 1650 36177
rect 1684 36143 1718 36177
rect 1752 36143 1786 36177
rect 1820 36143 1854 36177
rect 1888 36143 1922 36177
rect 1956 36143 1990 36177
rect 2024 36143 2058 36177
rect 2092 36143 2126 36177
rect 2160 36143 2194 36177
rect 2228 36143 2262 36177
rect 2296 36143 2330 36177
rect 2364 36143 2398 36177
rect 2432 36143 2466 36177
rect 2500 36143 2534 36177
rect 2568 36143 2602 36177
rect 2636 36143 2670 36177
rect 2704 36143 2738 36177
rect 2772 36143 2806 36177
rect 2840 36143 2874 36177
rect 2908 36143 2942 36177
rect 2976 36143 3010 36177
rect 3044 36143 3078 36177
rect 3112 36143 3146 36177
rect 3180 36143 3214 36177
rect 3248 36143 3282 36177
rect 3316 36143 3350 36177
rect 3384 36143 3418 36177
rect 3452 36143 3486 36177
rect 3520 36143 3554 36177
rect 3588 36143 3622 36177
rect 3656 36143 3690 36177
rect 3724 36143 3758 36177
rect 3792 36143 3826 36177
rect 3860 36143 3894 36177
rect 3928 36143 3962 36177
rect 3996 36143 4030 36177
rect 4064 36143 4098 36177
rect 4132 36143 4166 36177
rect 4200 36143 4234 36177
rect 4268 36143 4302 36177
rect 4336 36143 4370 36177
rect 4404 36143 4438 36177
rect 4472 36143 4506 36177
rect 4540 36143 4574 36177
rect 4608 36143 4642 36177
rect 4676 36143 4710 36177
rect 4744 36143 4778 36177
rect 4812 36143 4846 36177
rect 4880 36143 4914 36177
rect 4948 36143 4982 36177
rect 5016 36143 5050 36177
rect 5084 36143 5118 36177
rect 5152 36143 5186 36177
rect 5220 36143 5254 36177
rect 5288 36143 5322 36177
rect 5356 36143 5390 36177
rect 5424 36143 5458 36177
rect 5492 36143 5526 36177
rect 5560 36143 5594 36177
rect 5628 36143 5662 36177
rect 5696 36143 5730 36177
rect 5764 36143 5798 36177
rect 5832 36143 5866 36177
rect 5900 36143 5934 36177
rect 5968 36143 6002 36177
rect 6036 36143 6070 36177
rect 6104 36143 6138 36177
rect 6172 36143 6206 36177
rect 6240 36143 6274 36177
rect 6308 36143 6342 36177
rect 6376 36143 6410 36177
rect 6444 36143 6478 36177
rect 6512 36143 6546 36177
rect 6580 36143 6614 36177
rect 6648 36143 6682 36177
rect 6716 36143 6750 36177
rect 6784 36143 6818 36177
rect 6852 36143 6886 36177
rect 6920 36143 6954 36177
rect 6988 36143 7022 36177
rect 7056 36143 7090 36177
rect 7124 36143 7158 36177
rect 7192 36143 7226 36177
rect 7260 36143 7294 36177
rect 7328 36143 7362 36177
rect 7396 36143 7430 36177
rect 7464 36143 7498 36177
rect 7532 36143 7566 36177
rect 7600 36143 7634 36177
rect 7668 36143 7702 36177
rect 7736 36143 7770 36177
rect 7804 36143 7838 36177
rect 7872 36143 7906 36177
rect 7940 36143 7974 36177
rect 8008 36143 8042 36177
rect 8076 36143 8110 36177
rect 8144 36143 8178 36177
rect 8212 36143 8246 36177
rect 8280 36143 8314 36177
rect 8348 36143 8382 36177
rect 8416 36143 8450 36177
rect 8484 36143 8518 36177
rect 8552 36143 8586 36177
rect 8620 36143 8654 36177
rect 8688 36143 8722 36177
rect 8756 36143 8790 36177
rect 8824 36143 8858 36177
rect 8892 36143 8926 36177
rect 8960 36143 8994 36177
rect 9028 36143 9062 36177
rect 9096 36143 9130 36177
rect 9164 36143 9198 36177
rect 9232 36143 9266 36177
rect 9300 36143 9334 36177
rect 9368 36143 9402 36177
rect 9436 36143 9470 36177
rect 9504 36143 9538 36177
rect 9572 36143 9606 36177
rect 9640 36143 9674 36177
rect 9708 36143 9742 36177
rect 9776 36143 9810 36177
rect 9844 36143 9878 36177
rect 9912 36143 9946 36177
rect 9980 36143 10014 36177
rect 10048 36143 10082 36177
rect 10116 36143 10150 36177
rect 10184 36143 10218 36177
rect 10252 36143 10286 36177
rect 10320 36143 10354 36177
rect 10388 36143 10422 36177
rect 10456 36143 10490 36177
rect 10524 36143 10558 36177
rect 10592 36143 10626 36177
rect 10660 36143 10694 36177
rect 10728 36143 10762 36177
rect 10796 36143 10830 36177
rect 10864 36143 10898 36177
rect 10932 36143 10966 36177
rect 11000 36143 11034 36177
rect 11068 36143 11102 36177
rect 11136 36143 11170 36177
rect 11204 36143 11238 36177
rect 11272 36143 11306 36177
rect 11340 36143 11374 36177
rect 11408 36143 11442 36177
rect 11476 36143 11510 36177
rect 11544 36143 11578 36177
rect 11612 36143 11646 36177
rect 11680 36143 11714 36177
rect 11748 36143 11782 36177
rect 11816 36143 11850 36177
rect 11884 36143 11918 36177
rect 11952 36143 11986 36177
rect 12020 36143 12054 36177
rect 12088 36143 12122 36177
rect 12156 36143 12190 36177
rect 12224 36143 12258 36177
rect 12292 36143 12326 36177
rect 12360 36143 12394 36177
rect 12428 36143 12462 36177
rect 12496 36143 12530 36177
rect 12564 36143 12598 36177
rect 12632 36143 12666 36177
rect 12700 36143 12734 36177
rect 12768 36143 12802 36177
rect 12836 36143 12870 36177
rect 12904 36143 12938 36177
rect 12972 36143 13006 36177
rect 13040 36143 13074 36177
rect 13108 36143 13142 36177
rect 13176 36143 13210 36177
rect 13244 36143 13278 36177
rect 13312 36143 13346 36177
rect 13380 36143 13414 36177
rect 13448 36143 13482 36177
rect 13516 36143 13550 36177
rect 13584 36143 13618 36177
rect 13652 36143 13686 36177
rect 13720 36143 13754 36177
rect 13788 36143 13822 36177
rect 13856 36143 13890 36177
rect 13924 36143 13958 36177
rect 13992 36143 14026 36177
rect 14060 36143 14094 36177
rect 14128 36143 14162 36177
rect 14196 36143 14381 36177
rect 583 36093 14381 36143
rect 583 36050 715 36093
rect 583 36016 632 36050
rect 666 36016 715 36050
rect 583 35982 715 36016
rect 583 35948 632 35982
rect 666 35948 715 35982
rect 583 35914 715 35948
rect 583 35880 632 35914
rect 666 35880 715 35914
rect 583 35846 715 35880
rect 583 35812 632 35846
rect 666 35812 715 35846
rect 583 35778 715 35812
rect 583 35744 632 35778
rect 666 35744 715 35778
rect 583 35710 715 35744
rect 583 35676 632 35710
rect 666 35676 715 35710
rect 583 35642 715 35676
rect 583 35608 632 35642
rect 666 35608 715 35642
rect 583 35574 715 35608
rect 583 35540 632 35574
rect 666 35540 715 35574
rect 583 35506 715 35540
rect 583 35472 632 35506
rect 666 35472 715 35506
rect 583 35438 715 35472
rect 583 35404 632 35438
rect 666 35404 715 35438
rect 583 35370 715 35404
rect 583 35336 632 35370
rect 666 35336 715 35370
rect 583 35302 715 35336
rect 583 35268 632 35302
rect 666 35268 715 35302
rect 583 35234 715 35268
rect 583 35200 632 35234
rect 666 35200 715 35234
rect 583 35166 715 35200
rect 583 35132 632 35166
rect 666 35132 715 35166
rect 583 35098 715 35132
rect 583 35064 632 35098
rect 666 35064 715 35098
rect 583 35030 715 35064
rect 583 34996 632 35030
rect 666 34996 715 35030
rect 583 34962 715 34996
rect 583 34928 632 34962
rect 666 34928 715 34962
rect 583 34894 715 34928
rect 583 34860 632 34894
rect 666 34860 715 34894
rect 583 34826 715 34860
rect 583 34792 632 34826
rect 666 34792 715 34826
rect 583 34758 715 34792
rect 583 34724 632 34758
rect 666 34724 715 34758
rect 583 34690 715 34724
rect 14247 36050 14381 36093
rect 14247 36016 14297 36050
rect 14331 36016 14381 36050
rect 14247 35982 14381 36016
rect 14247 35948 14297 35982
rect 14331 35948 14381 35982
rect 14247 35914 14381 35948
rect 14247 35880 14297 35914
rect 14331 35880 14381 35914
rect 14247 35846 14381 35880
rect 14247 35812 14297 35846
rect 14331 35812 14381 35846
rect 14247 35778 14381 35812
rect 14247 35744 14297 35778
rect 14331 35744 14381 35778
rect 14247 35710 14381 35744
rect 14247 35676 14297 35710
rect 14331 35676 14381 35710
rect 14247 35642 14381 35676
rect 14247 35608 14297 35642
rect 14331 35608 14381 35642
rect 14247 35574 14381 35608
rect 14247 35540 14297 35574
rect 14331 35540 14381 35574
rect 14247 35506 14381 35540
rect 14247 35472 14297 35506
rect 14331 35472 14381 35506
rect 14247 35438 14381 35472
rect 14247 35404 14297 35438
rect 14331 35404 14381 35438
rect 14247 35370 14381 35404
rect 14247 35336 14297 35370
rect 14331 35336 14381 35370
rect 14247 35302 14381 35336
rect 14247 35268 14297 35302
rect 14331 35268 14381 35302
rect 14247 35234 14381 35268
rect 14247 35200 14297 35234
rect 14331 35200 14381 35234
rect 14247 35166 14381 35200
rect 14247 35132 14297 35166
rect 14331 35132 14381 35166
rect 14247 35098 14381 35132
rect 14247 35064 14297 35098
rect 14331 35064 14381 35098
rect 14247 35030 14381 35064
rect 14247 34996 14297 35030
rect 14331 34996 14381 35030
rect 14247 34962 14381 34996
rect 14247 34928 14297 34962
rect 14331 34928 14381 34962
rect 14247 34894 14381 34928
rect 14247 34860 14297 34894
rect 14331 34860 14381 34894
rect 14247 34826 14381 34860
rect 14247 34792 14297 34826
rect 14331 34792 14381 34826
rect 14247 34758 14381 34792
rect 14247 34724 14297 34758
rect 14331 34724 14381 34758
rect 583 34656 632 34690
rect 666 34656 715 34690
rect 583 34622 715 34656
rect 583 34588 632 34622
rect 666 34588 715 34622
rect 583 34554 715 34588
rect 583 34520 632 34554
rect 666 34520 715 34554
rect 583 34486 715 34520
rect 583 34452 632 34486
rect 666 34452 715 34486
rect 583 34418 715 34452
rect 583 34384 632 34418
rect 666 34384 715 34418
rect 583 34350 715 34384
rect 583 34316 632 34350
rect 666 34316 715 34350
rect 583 34282 715 34316
rect 583 34248 632 34282
rect 666 34248 715 34282
rect 583 34214 715 34248
rect 583 34180 632 34214
rect 666 34180 715 34214
rect 583 34146 715 34180
rect 583 34112 632 34146
rect 666 34112 715 34146
rect 583 34078 715 34112
rect 583 34044 632 34078
rect 666 34044 715 34078
rect 583 34010 715 34044
rect 583 33976 632 34010
rect 666 33976 715 34010
rect 583 33942 715 33976
rect 583 33908 632 33942
rect 666 33908 715 33942
rect 583 33874 715 33908
rect 583 33840 632 33874
rect 666 33840 715 33874
rect 583 33806 715 33840
rect 583 33772 632 33806
rect 666 33772 715 33806
rect 583 33738 715 33772
rect 583 33704 632 33738
rect 666 33704 715 33738
rect 583 33670 715 33704
rect 583 33636 632 33670
rect 666 33636 715 33670
rect 583 33602 715 33636
rect 583 33568 632 33602
rect 666 33568 715 33602
rect 583 33534 715 33568
rect 583 33500 632 33534
rect 666 33500 715 33534
rect 583 33466 715 33500
rect 583 33432 632 33466
rect 666 33432 715 33466
rect 583 33398 715 33432
rect 583 33364 632 33398
rect 666 33364 715 33398
rect 583 33330 715 33364
rect 583 33296 632 33330
rect 666 33296 715 33330
rect 583 33262 715 33296
rect 583 33228 632 33262
rect 666 33228 715 33262
rect 583 33194 715 33228
rect 583 33160 632 33194
rect 666 33160 715 33194
rect 583 33126 715 33160
rect 583 33092 632 33126
rect 666 33092 715 33126
rect 583 33058 715 33092
rect 583 33024 632 33058
rect 666 33024 715 33058
rect 583 32990 715 33024
rect 583 32956 632 32990
rect 666 32956 715 32990
rect 583 32922 715 32956
rect 583 32888 632 32922
rect 666 32888 715 32922
rect 583 32854 715 32888
rect 583 32820 632 32854
rect 666 32820 715 32854
rect 583 32786 715 32820
rect 583 32752 632 32786
rect 666 32752 715 32786
rect 583 32718 715 32752
rect 583 32684 632 32718
rect 666 32684 715 32718
rect 583 32650 715 32684
rect 583 32616 632 32650
rect 666 32616 715 32650
rect 583 32582 715 32616
rect 583 32548 632 32582
rect 666 32548 715 32582
rect 583 32514 715 32548
rect 583 32480 632 32514
rect 666 32480 715 32514
rect 583 32446 715 32480
rect 583 32412 632 32446
rect 666 32412 715 32446
rect 583 32378 715 32412
rect 583 32344 632 32378
rect 666 32344 715 32378
rect 583 32310 715 32344
rect 583 32276 632 32310
rect 666 32276 715 32310
rect 583 32242 715 32276
rect 583 32208 632 32242
rect 666 32208 715 32242
rect 583 32174 715 32208
rect 583 32140 632 32174
rect 666 32140 715 32174
rect 583 32106 715 32140
rect 583 32072 632 32106
rect 666 32072 715 32106
rect 583 32038 715 32072
rect 583 32004 632 32038
rect 666 32004 715 32038
rect 583 31970 715 32004
rect 583 31936 632 31970
rect 666 31936 715 31970
rect 583 31902 715 31936
rect 583 31868 632 31902
rect 666 31868 715 31902
rect 583 31834 715 31868
rect 583 31800 632 31834
rect 666 31800 715 31834
rect 583 31766 715 31800
rect 583 31732 632 31766
rect 666 31732 715 31766
rect 583 31698 715 31732
rect 583 31664 632 31698
rect 666 31664 715 31698
rect 583 31630 715 31664
rect 583 31596 632 31630
rect 666 31596 715 31630
rect 583 31562 715 31596
rect 583 31528 632 31562
rect 666 31528 715 31562
rect 583 31494 715 31528
rect 583 31460 632 31494
rect 666 31460 715 31494
rect 583 31426 715 31460
rect 583 31392 632 31426
rect 666 31392 715 31426
rect 583 31358 715 31392
rect 583 31324 632 31358
rect 666 31324 715 31358
rect 583 31290 715 31324
rect 583 31256 632 31290
rect 666 31256 715 31290
rect 583 31222 715 31256
rect 583 31188 632 31222
rect 666 31188 715 31222
rect 583 31154 715 31188
rect 583 31120 632 31154
rect 666 31120 715 31154
rect 583 31086 715 31120
rect 583 31052 632 31086
rect 666 31052 715 31086
rect 583 31018 715 31052
rect 583 30984 632 31018
rect 666 30984 715 31018
rect 583 30950 715 30984
rect 583 30916 632 30950
rect 666 30916 715 30950
rect 583 30882 715 30916
rect 583 30848 632 30882
rect 666 30848 715 30882
rect 583 30814 715 30848
rect 583 30780 632 30814
rect 666 30780 715 30814
rect 583 30746 715 30780
rect 583 30712 632 30746
rect 666 30712 715 30746
rect 583 30678 715 30712
rect 583 30644 632 30678
rect 666 30644 715 30678
rect 583 30610 715 30644
rect 583 30576 632 30610
rect 666 30576 715 30610
rect 583 30542 715 30576
rect 583 30508 632 30542
rect 666 30508 715 30542
rect 583 30474 715 30508
rect 583 30440 632 30474
rect 666 30440 715 30474
rect 583 30406 715 30440
rect 583 30372 632 30406
rect 666 30372 715 30406
rect 583 30338 715 30372
rect 583 30304 632 30338
rect 666 30304 715 30338
rect 583 30270 715 30304
rect 583 30236 632 30270
rect 666 30236 715 30270
rect 583 30202 715 30236
rect 583 30168 632 30202
rect 666 30168 715 30202
rect 583 30134 715 30168
rect 583 30100 632 30134
rect 666 30100 715 30134
rect 583 30066 715 30100
rect 583 30032 632 30066
rect 666 30032 715 30066
rect 583 29998 715 30032
rect 583 29964 632 29998
rect 666 29964 715 29998
rect 583 29930 715 29964
rect 583 29896 632 29930
rect 666 29896 715 29930
rect 583 29862 715 29896
rect 583 29828 632 29862
rect 666 29828 715 29862
rect 583 29794 715 29828
rect 583 29760 632 29794
rect 666 29760 715 29794
rect 583 29726 715 29760
rect 583 29692 632 29726
rect 666 29692 715 29726
rect 583 29658 715 29692
rect 583 29624 632 29658
rect 666 29624 715 29658
rect 583 29590 715 29624
rect 583 29556 632 29590
rect 666 29556 715 29590
rect 583 29522 715 29556
rect 583 29488 632 29522
rect 666 29488 715 29522
rect 583 29454 715 29488
rect 583 29420 632 29454
rect 666 29420 715 29454
rect 583 29386 715 29420
rect 583 29352 632 29386
rect 666 29352 715 29386
rect 583 29318 715 29352
rect 583 29284 632 29318
rect 666 29284 715 29318
rect 583 29250 715 29284
rect 583 29216 632 29250
rect 666 29216 715 29250
rect 583 29182 715 29216
rect 583 29148 632 29182
rect 666 29148 715 29182
rect 583 29114 715 29148
rect 583 29080 632 29114
rect 666 29080 715 29114
rect 583 29046 715 29080
rect 583 29012 632 29046
rect 666 29012 715 29046
rect 583 28978 715 29012
rect 583 28944 632 28978
rect 666 28944 715 28978
rect 583 28910 715 28944
rect 583 28876 632 28910
rect 666 28876 715 28910
rect 583 28842 715 28876
rect 583 28808 632 28842
rect 666 28808 715 28842
rect 583 28774 715 28808
rect 583 28740 632 28774
rect 666 28740 715 28774
rect 583 28706 715 28740
rect 583 28672 632 28706
rect 666 28672 715 28706
rect 583 28638 715 28672
rect 583 28604 632 28638
rect 666 28604 715 28638
rect 583 28570 715 28604
rect 583 28536 632 28570
rect 666 28536 715 28570
rect 583 28502 715 28536
rect 583 28468 632 28502
rect 666 28468 715 28502
rect 583 28434 715 28468
rect 583 28400 632 28434
rect 666 28400 715 28434
rect 583 28366 715 28400
rect 583 28332 632 28366
rect 666 28332 715 28366
rect 583 28298 715 28332
rect 583 28264 632 28298
rect 666 28264 715 28298
rect 583 28230 715 28264
rect 583 28196 632 28230
rect 666 28196 715 28230
rect 583 28162 715 28196
rect 583 28128 632 28162
rect 666 28128 715 28162
rect 583 28094 715 28128
rect 583 28060 632 28094
rect 666 28060 715 28094
rect 583 28026 715 28060
rect 583 27992 632 28026
rect 666 27992 715 28026
rect 583 27958 715 27992
rect 583 27924 632 27958
rect 666 27924 715 27958
rect 583 27890 715 27924
rect 583 27856 632 27890
rect 666 27856 715 27890
rect 583 27822 715 27856
rect 583 27788 632 27822
rect 666 27788 715 27822
rect 583 27754 715 27788
rect 583 27720 632 27754
rect 666 27720 715 27754
rect 583 27686 715 27720
rect 583 27652 632 27686
rect 666 27652 715 27686
rect 583 27618 715 27652
rect 583 27584 632 27618
rect 666 27584 715 27618
rect 583 27550 715 27584
rect 583 27516 632 27550
rect 666 27516 715 27550
rect 583 27482 715 27516
rect 583 27448 632 27482
rect 666 27448 715 27482
rect 583 27414 715 27448
rect 583 27380 632 27414
rect 666 27380 715 27414
rect 583 27346 715 27380
rect 583 27312 632 27346
rect 666 27312 715 27346
rect 583 27278 715 27312
rect 583 27244 632 27278
rect 666 27244 715 27278
rect 583 27210 715 27244
rect 583 27176 632 27210
rect 666 27176 715 27210
rect 583 27142 715 27176
rect 583 27108 632 27142
rect 666 27108 715 27142
rect 583 27074 715 27108
rect 583 27040 632 27074
rect 666 27040 715 27074
rect 583 27006 715 27040
rect 583 26972 632 27006
rect 666 26972 715 27006
rect 583 26938 715 26972
rect 583 26904 632 26938
rect 666 26904 715 26938
rect 583 26870 715 26904
rect 583 26836 632 26870
rect 666 26836 715 26870
rect 583 26802 715 26836
rect 583 26768 632 26802
rect 666 26768 715 26802
rect 583 26734 715 26768
rect 583 26700 632 26734
rect 666 26700 715 26734
rect 583 26666 715 26700
rect 583 26632 632 26666
rect 666 26632 715 26666
rect 583 26598 715 26632
rect 583 26564 632 26598
rect 666 26564 715 26598
rect 583 26530 715 26564
rect 583 26496 632 26530
rect 666 26496 715 26530
rect 583 26462 715 26496
rect 583 26428 632 26462
rect 666 26428 715 26462
rect 583 26394 715 26428
rect 583 26360 632 26394
rect 666 26360 715 26394
rect 583 26326 715 26360
rect 583 26292 632 26326
rect 666 26292 715 26326
rect 583 26258 715 26292
rect 583 26224 632 26258
rect 666 26224 715 26258
rect 583 26190 715 26224
rect 583 26156 632 26190
rect 666 26156 715 26190
rect 583 26122 715 26156
rect 583 26088 632 26122
rect 666 26088 715 26122
rect 583 26054 715 26088
rect 583 26020 632 26054
rect 666 26020 715 26054
rect 583 25986 715 26020
rect 583 25952 632 25986
rect 666 25952 715 25986
rect 583 25918 715 25952
rect 583 25884 632 25918
rect 666 25884 715 25918
rect 583 25850 715 25884
rect 583 25816 632 25850
rect 666 25816 715 25850
rect 583 25782 715 25816
rect 583 25748 632 25782
rect 666 25748 715 25782
rect 583 25714 715 25748
rect 583 25680 632 25714
rect 666 25680 715 25714
rect 583 25646 715 25680
rect 583 25612 632 25646
rect 666 25612 715 25646
rect 583 25578 715 25612
rect 583 25544 632 25578
rect 666 25544 715 25578
rect 583 25510 715 25544
rect 583 25476 632 25510
rect 666 25476 715 25510
rect 583 25442 715 25476
rect 583 25408 632 25442
rect 666 25408 715 25442
rect 583 25374 715 25408
rect 583 25340 632 25374
rect 666 25340 715 25374
rect 583 25306 715 25340
rect 583 25272 632 25306
rect 666 25272 715 25306
rect 583 25238 715 25272
rect 583 25204 632 25238
rect 666 25204 715 25238
rect 583 25170 715 25204
rect 583 25136 632 25170
rect 666 25136 715 25170
rect 583 25102 715 25136
rect 583 25068 632 25102
rect 666 25068 715 25102
rect 583 25034 715 25068
rect 583 25000 632 25034
rect 666 25000 715 25034
rect 583 24966 715 25000
rect 583 24932 632 24966
rect 666 24932 715 24966
rect 583 24898 715 24932
rect 583 24864 632 24898
rect 666 24864 715 24898
rect 583 24830 715 24864
rect 583 24796 632 24830
rect 666 24796 715 24830
rect 583 24762 715 24796
rect 583 24728 632 24762
rect 666 24728 715 24762
rect 583 24694 715 24728
rect 583 24660 632 24694
rect 666 24660 715 24694
rect 583 24626 715 24660
rect 583 24592 632 24626
rect 666 24592 715 24626
rect 583 24558 715 24592
rect 583 24524 632 24558
rect 666 24524 715 24558
rect 583 24490 715 24524
rect 583 24456 632 24490
rect 666 24456 715 24490
rect 583 24422 715 24456
rect 583 24388 632 24422
rect 666 24388 715 24422
rect 583 24354 715 24388
rect 583 24320 632 24354
rect 666 24320 715 24354
rect 583 24286 715 24320
rect 583 24252 632 24286
rect 666 24252 715 24286
rect 583 24218 715 24252
rect 583 24184 632 24218
rect 666 24184 715 24218
rect 583 24150 715 24184
rect 583 24116 632 24150
rect 666 24116 715 24150
rect 583 24082 715 24116
rect 583 24048 632 24082
rect 666 24048 715 24082
rect 583 24014 715 24048
rect 583 23980 632 24014
rect 666 23980 715 24014
rect 583 23946 715 23980
rect 583 23912 632 23946
rect 666 23912 715 23946
rect 583 23878 715 23912
rect 583 23844 632 23878
rect 666 23844 715 23878
rect 583 23810 715 23844
rect 583 23776 632 23810
rect 666 23776 715 23810
rect 583 23742 715 23776
rect 583 23708 632 23742
rect 666 23708 715 23742
rect 583 23674 715 23708
rect 583 23640 632 23674
rect 666 23640 715 23674
rect 583 23606 715 23640
rect 583 23572 632 23606
rect 666 23572 715 23606
rect 583 23538 715 23572
rect 583 23504 632 23538
rect 666 23504 715 23538
rect 583 23470 715 23504
rect 583 23436 632 23470
rect 666 23436 715 23470
rect 583 23402 715 23436
rect 583 23368 632 23402
rect 666 23368 715 23402
rect 583 23334 715 23368
rect 583 23300 632 23334
rect 666 23300 715 23334
rect 583 23266 715 23300
rect 583 23232 632 23266
rect 666 23232 715 23266
rect 583 23198 715 23232
rect 583 23164 632 23198
rect 666 23164 715 23198
rect 583 23130 715 23164
rect 583 23096 632 23130
rect 666 23096 715 23130
rect 583 23062 715 23096
rect 583 23028 632 23062
rect 666 23028 715 23062
rect 583 22994 715 23028
rect 583 22960 632 22994
rect 666 22960 715 22994
rect 583 22926 715 22960
rect 583 22892 632 22926
rect 666 22892 715 22926
rect 583 22858 715 22892
rect 583 22824 632 22858
rect 666 22824 715 22858
rect 583 22790 715 22824
rect 583 22756 632 22790
rect 666 22756 715 22790
rect 583 22722 715 22756
rect 583 22688 632 22722
rect 666 22688 715 22722
rect 583 22654 715 22688
rect 583 22620 632 22654
rect 666 22620 715 22654
rect 583 22586 715 22620
rect 583 22552 632 22586
rect 666 22552 715 22586
rect 583 22518 715 22552
rect 583 22484 632 22518
rect 666 22484 715 22518
rect 583 22450 715 22484
rect 583 22416 632 22450
rect 666 22416 715 22450
rect 583 22382 715 22416
rect 583 22348 632 22382
rect 666 22348 715 22382
rect 583 22314 715 22348
rect 583 22280 632 22314
rect 666 22280 715 22314
rect 583 22246 715 22280
rect 583 22212 632 22246
rect 666 22212 715 22246
rect 583 22178 715 22212
rect 583 22144 632 22178
rect 666 22144 715 22178
rect 583 22110 715 22144
rect 583 22076 632 22110
rect 666 22076 715 22110
rect 583 22042 715 22076
rect 583 22008 632 22042
rect 666 22008 715 22042
rect 583 21974 715 22008
rect 583 21940 632 21974
rect 666 21940 715 21974
rect 583 21906 715 21940
rect 583 21872 632 21906
rect 666 21872 715 21906
rect 583 21838 715 21872
rect 583 21804 632 21838
rect 666 21804 715 21838
rect 583 21770 715 21804
rect 583 21736 632 21770
rect 666 21736 715 21770
rect 583 21702 715 21736
rect 583 21668 632 21702
rect 666 21668 715 21702
rect 583 21634 715 21668
rect 583 21600 632 21634
rect 666 21600 715 21634
rect 583 21566 715 21600
rect 583 21532 632 21566
rect 666 21532 715 21566
rect 583 21498 715 21532
rect 583 21464 632 21498
rect 666 21464 715 21498
rect 583 21430 715 21464
rect 583 21396 632 21430
rect 666 21396 715 21430
rect 583 21362 715 21396
rect 583 21328 632 21362
rect 666 21328 715 21362
rect 583 21294 715 21328
rect 583 21260 632 21294
rect 666 21260 715 21294
rect 583 21226 715 21260
rect 583 21192 632 21226
rect 666 21192 715 21226
rect 583 21158 715 21192
rect 583 21124 632 21158
rect 666 21124 715 21158
rect 583 21090 715 21124
rect 583 21056 632 21090
rect 666 21056 715 21090
rect 583 21022 715 21056
rect 583 20988 632 21022
rect 666 20988 715 21022
rect 583 20954 715 20988
rect 583 20920 632 20954
rect 666 20920 715 20954
rect 583 20886 715 20920
rect 583 20852 632 20886
rect 666 20852 715 20886
rect 583 20818 715 20852
rect 583 20784 632 20818
rect 666 20784 715 20818
rect 583 20750 715 20784
rect 583 20716 632 20750
rect 666 20716 715 20750
rect 583 20682 715 20716
rect 583 20648 632 20682
rect 666 20648 715 20682
rect 583 20614 715 20648
rect 583 20580 632 20614
rect 666 20580 715 20614
rect 583 20546 715 20580
rect 583 20512 632 20546
rect 666 20512 715 20546
rect 583 20478 715 20512
rect 583 20444 632 20478
rect 666 20444 715 20478
rect 583 20410 715 20444
rect 583 20376 632 20410
rect 666 20376 715 20410
rect 583 20342 715 20376
rect 583 20308 632 20342
rect 666 20308 715 20342
rect 583 20274 715 20308
rect 583 20240 632 20274
rect 666 20240 715 20274
rect 583 20206 715 20240
rect 583 20172 632 20206
rect 666 20172 715 20206
rect 583 20138 715 20172
rect 583 20104 632 20138
rect 666 20104 715 20138
rect 583 20070 715 20104
rect 583 20036 632 20070
rect 666 20036 715 20070
rect 583 20002 715 20036
rect 583 19968 632 20002
rect 666 19968 715 20002
rect 583 19934 715 19968
rect 583 19900 632 19934
rect 666 19900 715 19934
rect 583 19866 715 19900
rect 583 19832 632 19866
rect 666 19832 715 19866
rect 583 19798 715 19832
rect 583 19764 632 19798
rect 666 19764 715 19798
rect 583 19730 715 19764
rect 583 19696 632 19730
rect 666 19696 715 19730
rect 583 19662 715 19696
rect 583 19628 632 19662
rect 666 19628 715 19662
rect 583 19594 715 19628
rect 583 19560 632 19594
rect 666 19560 715 19594
rect 583 19526 715 19560
rect 583 19492 632 19526
rect 666 19492 715 19526
rect 583 19458 715 19492
rect 583 19424 632 19458
rect 666 19424 715 19458
rect 583 19390 715 19424
rect 583 19356 632 19390
rect 666 19356 715 19390
rect 583 19322 715 19356
rect 583 19288 632 19322
rect 666 19288 715 19322
rect 583 19254 715 19288
rect 583 19220 632 19254
rect 666 19220 715 19254
rect 583 19186 715 19220
rect 583 19152 632 19186
rect 666 19152 715 19186
rect 583 19118 715 19152
rect 583 19084 632 19118
rect 666 19084 715 19118
rect 583 19050 715 19084
rect 583 19016 632 19050
rect 666 19016 715 19050
rect 583 18982 715 19016
rect 583 18948 632 18982
rect 666 18948 715 18982
rect 583 18914 715 18948
rect 583 18880 632 18914
rect 666 18880 715 18914
rect 583 18846 715 18880
rect 583 18812 632 18846
rect 666 18812 715 18846
rect 583 18778 715 18812
rect 583 18744 632 18778
rect 666 18744 715 18778
rect 583 18710 715 18744
rect 583 18676 632 18710
rect 666 18676 715 18710
rect 583 18642 715 18676
rect 583 18608 632 18642
rect 666 18608 715 18642
rect 583 18574 715 18608
rect 583 18540 632 18574
rect 666 18540 715 18574
rect 583 18506 715 18540
rect 583 18472 632 18506
rect 666 18472 715 18506
rect 583 18438 715 18472
rect 583 18404 632 18438
rect 666 18404 715 18438
rect 583 18370 715 18404
rect 583 18336 632 18370
rect 666 18336 715 18370
rect 583 18302 715 18336
rect 583 18268 632 18302
rect 666 18268 715 18302
rect 583 18234 715 18268
rect 583 18200 632 18234
rect 666 18200 715 18234
rect 583 18166 715 18200
rect 583 18132 632 18166
rect 666 18132 715 18166
rect 583 18098 715 18132
rect 583 18064 632 18098
rect 666 18064 715 18098
rect 583 18030 715 18064
rect 583 17996 632 18030
rect 666 17996 715 18030
rect 583 17962 715 17996
rect 583 17928 632 17962
rect 666 17928 715 17962
rect 583 17894 715 17928
rect 583 17860 632 17894
rect 666 17860 715 17894
rect 583 17826 715 17860
rect 583 17792 632 17826
rect 666 17792 715 17826
rect 583 17758 715 17792
rect 583 17724 632 17758
rect 666 17724 715 17758
rect 583 17690 715 17724
rect 583 17656 632 17690
rect 666 17656 715 17690
rect 583 17622 715 17656
rect 583 17588 632 17622
rect 666 17588 715 17622
rect 583 17554 715 17588
rect 583 17520 632 17554
rect 666 17520 715 17554
rect 583 17486 715 17520
rect 583 17452 632 17486
rect 666 17452 715 17486
rect 583 17418 715 17452
rect 583 17384 632 17418
rect 666 17384 715 17418
rect 583 17350 715 17384
rect 583 17316 632 17350
rect 666 17316 715 17350
rect 583 17282 715 17316
rect 583 17248 632 17282
rect 666 17248 715 17282
rect 583 17214 715 17248
rect 583 17180 632 17214
rect 666 17180 715 17214
rect 583 17146 715 17180
rect 583 17112 632 17146
rect 666 17112 715 17146
rect 583 17078 715 17112
rect 583 17044 632 17078
rect 666 17044 715 17078
rect 583 17010 715 17044
rect 583 16976 632 17010
rect 666 16976 715 17010
rect 583 16942 715 16976
rect 583 16908 632 16942
rect 666 16908 715 16942
rect 583 16874 715 16908
rect 583 16840 632 16874
rect 666 16840 715 16874
rect 583 16806 715 16840
rect 583 16772 632 16806
rect 666 16772 715 16806
rect 583 16738 715 16772
rect 583 16704 632 16738
rect 666 16704 715 16738
rect 583 16670 715 16704
rect 583 16636 632 16670
rect 666 16636 715 16670
rect 583 16602 715 16636
rect 583 16568 632 16602
rect 666 16568 715 16602
rect 583 16534 715 16568
rect 583 16500 632 16534
rect 666 16500 715 16534
rect 583 16466 715 16500
rect 583 16432 632 16466
rect 666 16432 715 16466
rect 583 16398 715 16432
rect 583 16364 632 16398
rect 666 16364 715 16398
rect 583 16330 715 16364
rect 583 16296 632 16330
rect 666 16296 715 16330
rect 583 16262 715 16296
rect 583 16228 632 16262
rect 666 16228 715 16262
rect 583 16194 715 16228
rect 583 16160 632 16194
rect 666 16160 715 16194
rect 583 16126 715 16160
rect 583 16092 632 16126
rect 666 16092 715 16126
rect 583 16058 715 16092
rect 583 16024 632 16058
rect 666 16024 715 16058
rect 583 15990 715 16024
rect 583 15956 632 15990
rect 666 15956 715 15990
rect 583 15922 715 15956
rect 583 15888 632 15922
rect 666 15888 715 15922
rect 583 15854 715 15888
rect 583 15820 632 15854
rect 666 15820 715 15854
rect 583 15786 715 15820
rect 583 15752 632 15786
rect 666 15752 715 15786
rect 583 15718 715 15752
rect 583 15684 632 15718
rect 666 15684 715 15718
rect 583 15650 715 15684
rect 583 15616 632 15650
rect 666 15616 715 15650
rect 583 15582 715 15616
rect 583 15548 632 15582
rect 666 15548 715 15582
rect 583 15514 715 15548
rect 583 15480 632 15514
rect 666 15480 715 15514
rect 583 15446 715 15480
rect 583 15412 632 15446
rect 666 15412 715 15446
rect 583 15378 715 15412
rect 583 15344 632 15378
rect 666 15344 715 15378
rect 583 15310 715 15344
rect 583 15276 632 15310
rect 666 15276 715 15310
rect 583 15242 715 15276
rect 583 15208 632 15242
rect 666 15208 715 15242
rect 583 15174 715 15208
rect 1659 28879 13357 28909
rect 1659 28505 2119 28879
rect 12897 28505 13357 28879
rect 1659 28475 13357 28505
rect 1659 28422 2093 28475
rect 1659 27504 1689 28422
rect 2063 27504 2093 28422
rect 1659 27451 2093 27504
rect 12923 28422 13357 28475
rect 12923 27504 12953 28422
rect 13327 27504 13357 28422
rect 12923 27451 13357 27504
rect 1659 27421 13357 27451
rect 1659 27047 2119 27421
rect 12897 27047 13357 27421
rect 1659 27017 13357 27047
rect 14247 34690 14381 34724
rect 14247 34656 14297 34690
rect 14331 34656 14381 34690
rect 14247 34622 14381 34656
rect 14247 34588 14297 34622
rect 14331 34588 14381 34622
rect 14247 34554 14381 34588
rect 14247 34520 14297 34554
rect 14331 34520 14381 34554
rect 14247 34486 14381 34520
rect 14247 34452 14297 34486
rect 14331 34452 14381 34486
rect 14247 34418 14381 34452
rect 14247 34384 14297 34418
rect 14331 34384 14381 34418
rect 14247 34350 14381 34384
rect 14247 34316 14297 34350
rect 14331 34316 14381 34350
rect 14247 34282 14381 34316
rect 14247 34248 14297 34282
rect 14331 34248 14381 34282
rect 14247 34214 14381 34248
rect 14247 34180 14297 34214
rect 14331 34180 14381 34214
rect 14247 34146 14381 34180
rect 14247 34112 14297 34146
rect 14331 34112 14381 34146
rect 14247 34078 14381 34112
rect 14247 34044 14297 34078
rect 14331 34044 14381 34078
rect 14247 34010 14381 34044
rect 14247 33976 14297 34010
rect 14331 33976 14381 34010
rect 14247 33942 14381 33976
rect 14247 33908 14297 33942
rect 14331 33908 14381 33942
rect 14247 33874 14381 33908
rect 14247 33840 14297 33874
rect 14331 33840 14381 33874
rect 14247 33806 14381 33840
rect 14247 33772 14297 33806
rect 14331 33772 14381 33806
rect 14247 33738 14381 33772
rect 14247 33704 14297 33738
rect 14331 33704 14381 33738
rect 14247 33670 14381 33704
rect 14247 33636 14297 33670
rect 14331 33636 14381 33670
rect 14247 33602 14381 33636
rect 14247 33568 14297 33602
rect 14331 33568 14381 33602
rect 14247 33534 14381 33568
rect 14247 33500 14297 33534
rect 14331 33500 14381 33534
rect 14247 33466 14381 33500
rect 14247 33432 14297 33466
rect 14331 33432 14381 33466
rect 14247 33398 14381 33432
rect 14247 33364 14297 33398
rect 14331 33364 14381 33398
rect 14247 33330 14381 33364
rect 14247 33296 14297 33330
rect 14331 33296 14381 33330
rect 14247 33262 14381 33296
rect 14247 33228 14297 33262
rect 14331 33228 14381 33262
rect 14247 33194 14381 33228
rect 14247 33160 14297 33194
rect 14331 33160 14381 33194
rect 14247 33126 14381 33160
rect 14247 33092 14297 33126
rect 14331 33092 14381 33126
rect 14247 33058 14381 33092
rect 14247 33024 14297 33058
rect 14331 33024 14381 33058
rect 14247 32990 14381 33024
rect 14247 32956 14297 32990
rect 14331 32956 14381 32990
rect 14247 32922 14381 32956
rect 14247 32888 14297 32922
rect 14331 32888 14381 32922
rect 14247 32854 14381 32888
rect 14247 32820 14297 32854
rect 14331 32820 14381 32854
rect 14247 32786 14381 32820
rect 14247 32752 14297 32786
rect 14331 32752 14381 32786
rect 14247 32718 14381 32752
rect 14247 32684 14297 32718
rect 14331 32684 14381 32718
rect 14247 32650 14381 32684
rect 14247 32616 14297 32650
rect 14331 32616 14381 32650
rect 14247 32582 14381 32616
rect 14247 32548 14297 32582
rect 14331 32548 14381 32582
rect 14247 32514 14381 32548
rect 14247 32480 14297 32514
rect 14331 32480 14381 32514
rect 14247 32446 14381 32480
rect 14247 32412 14297 32446
rect 14331 32412 14381 32446
rect 14247 32378 14381 32412
rect 14247 32344 14297 32378
rect 14331 32344 14381 32378
rect 14247 32310 14381 32344
rect 14247 32276 14297 32310
rect 14331 32276 14381 32310
rect 14247 32242 14381 32276
rect 14247 32208 14297 32242
rect 14331 32208 14381 32242
rect 14247 32174 14381 32208
rect 14247 32140 14297 32174
rect 14331 32140 14381 32174
rect 14247 32106 14381 32140
rect 14247 32072 14297 32106
rect 14331 32072 14381 32106
rect 14247 32038 14381 32072
rect 14247 32004 14297 32038
rect 14331 32004 14381 32038
rect 14247 31970 14381 32004
rect 14247 31936 14297 31970
rect 14331 31936 14381 31970
rect 14247 31902 14381 31936
rect 14247 31868 14297 31902
rect 14331 31868 14381 31902
rect 14247 31834 14381 31868
rect 14247 31800 14297 31834
rect 14331 31800 14381 31834
rect 14247 31766 14381 31800
rect 14247 31732 14297 31766
rect 14331 31732 14381 31766
rect 14247 31698 14381 31732
rect 14247 31664 14297 31698
rect 14331 31664 14381 31698
rect 14247 31630 14381 31664
rect 14247 31596 14297 31630
rect 14331 31596 14381 31630
rect 14247 31562 14381 31596
rect 14247 31528 14297 31562
rect 14331 31528 14381 31562
rect 14247 31494 14381 31528
rect 14247 31460 14297 31494
rect 14331 31460 14381 31494
rect 14247 31426 14381 31460
rect 14247 31392 14297 31426
rect 14331 31392 14381 31426
rect 14247 31358 14381 31392
rect 14247 31324 14297 31358
rect 14331 31324 14381 31358
rect 14247 31290 14381 31324
rect 14247 31256 14297 31290
rect 14331 31256 14381 31290
rect 14247 31222 14381 31256
rect 14247 31188 14297 31222
rect 14331 31188 14381 31222
rect 14247 31154 14381 31188
rect 14247 31120 14297 31154
rect 14331 31120 14381 31154
rect 14247 31086 14381 31120
rect 14247 31052 14297 31086
rect 14331 31052 14381 31086
rect 14247 31018 14381 31052
rect 14247 30984 14297 31018
rect 14331 30984 14381 31018
rect 14247 30950 14381 30984
rect 14247 30916 14297 30950
rect 14331 30916 14381 30950
rect 14247 30882 14381 30916
rect 14247 30848 14297 30882
rect 14331 30848 14381 30882
rect 14247 30814 14381 30848
rect 14247 30780 14297 30814
rect 14331 30780 14381 30814
rect 14247 30746 14381 30780
rect 14247 30712 14297 30746
rect 14331 30712 14381 30746
rect 14247 30678 14381 30712
rect 14247 30644 14297 30678
rect 14331 30644 14381 30678
rect 14247 30610 14381 30644
rect 14247 30576 14297 30610
rect 14331 30576 14381 30610
rect 14247 30542 14381 30576
rect 14247 30508 14297 30542
rect 14331 30508 14381 30542
rect 14247 30474 14381 30508
rect 14247 30440 14297 30474
rect 14331 30440 14381 30474
rect 14247 30406 14381 30440
rect 14247 30372 14297 30406
rect 14331 30372 14381 30406
rect 14247 30338 14381 30372
rect 14247 30304 14297 30338
rect 14331 30304 14381 30338
rect 14247 30270 14381 30304
rect 14247 30236 14297 30270
rect 14331 30236 14381 30270
rect 14247 30202 14381 30236
rect 14247 30168 14297 30202
rect 14331 30168 14381 30202
rect 14247 30134 14381 30168
rect 14247 30100 14297 30134
rect 14331 30100 14381 30134
rect 14247 30066 14381 30100
rect 14247 30032 14297 30066
rect 14331 30032 14381 30066
rect 14247 29998 14381 30032
rect 14247 29964 14297 29998
rect 14331 29964 14381 29998
rect 14247 29930 14381 29964
rect 14247 29896 14297 29930
rect 14331 29896 14381 29930
rect 14247 29862 14381 29896
rect 14247 29828 14297 29862
rect 14331 29828 14381 29862
rect 14247 29794 14381 29828
rect 14247 29760 14297 29794
rect 14331 29760 14381 29794
rect 14247 29726 14381 29760
rect 14247 29692 14297 29726
rect 14331 29692 14381 29726
rect 14247 29658 14381 29692
rect 14247 29624 14297 29658
rect 14331 29624 14381 29658
rect 14247 29590 14381 29624
rect 14247 29556 14297 29590
rect 14331 29556 14381 29590
rect 14247 29522 14381 29556
rect 14247 29488 14297 29522
rect 14331 29488 14381 29522
rect 14247 29454 14381 29488
rect 14247 29420 14297 29454
rect 14331 29420 14381 29454
rect 14247 29386 14381 29420
rect 14247 29352 14297 29386
rect 14331 29352 14381 29386
rect 14247 29318 14381 29352
rect 14247 29284 14297 29318
rect 14331 29284 14381 29318
rect 14247 29250 14381 29284
rect 14247 29216 14297 29250
rect 14331 29216 14381 29250
rect 14247 29182 14381 29216
rect 14247 29148 14297 29182
rect 14331 29148 14381 29182
rect 14247 29114 14381 29148
rect 14247 29080 14297 29114
rect 14331 29080 14381 29114
rect 14247 29046 14381 29080
rect 14247 29012 14297 29046
rect 14331 29012 14381 29046
rect 14247 28978 14381 29012
rect 14247 28944 14297 28978
rect 14331 28944 14381 28978
rect 14247 28910 14381 28944
rect 14247 28876 14297 28910
rect 14331 28876 14381 28910
rect 14247 28842 14381 28876
rect 14247 28808 14297 28842
rect 14331 28808 14381 28842
rect 14247 28774 14381 28808
rect 14247 28740 14297 28774
rect 14331 28740 14381 28774
rect 14247 28706 14381 28740
rect 14247 28672 14297 28706
rect 14331 28672 14381 28706
rect 14247 28638 14381 28672
rect 14247 28604 14297 28638
rect 14331 28604 14381 28638
rect 14247 28570 14381 28604
rect 14247 28536 14297 28570
rect 14331 28536 14381 28570
rect 14247 28502 14381 28536
rect 14247 28468 14297 28502
rect 14331 28468 14381 28502
rect 14247 28434 14381 28468
rect 14247 28400 14297 28434
rect 14331 28400 14381 28434
rect 14247 28366 14381 28400
rect 14247 28332 14297 28366
rect 14331 28332 14381 28366
rect 14247 28298 14381 28332
rect 14247 28264 14297 28298
rect 14331 28264 14381 28298
rect 14247 28230 14381 28264
rect 14247 28196 14297 28230
rect 14331 28196 14381 28230
rect 14247 28162 14381 28196
rect 14247 28128 14297 28162
rect 14331 28128 14381 28162
rect 14247 28094 14381 28128
rect 14247 28060 14297 28094
rect 14331 28060 14381 28094
rect 14247 28026 14381 28060
rect 14247 27992 14297 28026
rect 14331 27992 14381 28026
rect 14247 27958 14381 27992
rect 14247 27924 14297 27958
rect 14331 27924 14381 27958
rect 14247 27890 14381 27924
rect 14247 27856 14297 27890
rect 14331 27856 14381 27890
rect 14247 27822 14381 27856
rect 14247 27788 14297 27822
rect 14331 27788 14381 27822
rect 14247 27754 14381 27788
rect 14247 27720 14297 27754
rect 14331 27720 14381 27754
rect 14247 27686 14381 27720
rect 14247 27652 14297 27686
rect 14331 27652 14381 27686
rect 14247 27618 14381 27652
rect 14247 27584 14297 27618
rect 14331 27584 14381 27618
rect 14247 27550 14381 27584
rect 14247 27516 14297 27550
rect 14331 27516 14381 27550
rect 14247 27482 14381 27516
rect 14247 27448 14297 27482
rect 14331 27448 14381 27482
rect 14247 27414 14381 27448
rect 14247 27380 14297 27414
rect 14331 27380 14381 27414
rect 14247 27346 14381 27380
rect 14247 27312 14297 27346
rect 14331 27312 14381 27346
rect 14247 27278 14381 27312
rect 14247 27244 14297 27278
rect 14331 27244 14381 27278
rect 14247 27210 14381 27244
rect 14247 27176 14297 27210
rect 14331 27176 14381 27210
rect 14247 27142 14381 27176
rect 14247 27108 14297 27142
rect 14331 27108 14381 27142
rect 14247 27074 14381 27108
rect 14247 27040 14297 27074
rect 14331 27040 14381 27074
rect 14247 27006 14381 27040
rect 14247 26972 14297 27006
rect 14331 26972 14381 27006
rect 14247 26938 14381 26972
rect 14247 26904 14297 26938
rect 14331 26904 14381 26938
rect 14247 26870 14381 26904
rect 14247 26836 14297 26870
rect 14331 26836 14381 26870
rect 14247 26802 14381 26836
rect 14247 26768 14297 26802
rect 14331 26768 14381 26802
rect 14247 26734 14381 26768
rect 14247 26700 14297 26734
rect 14331 26700 14381 26734
rect 14247 26666 14381 26700
rect 14247 26632 14297 26666
rect 14331 26632 14381 26666
rect 14247 26598 14381 26632
rect 14247 26564 14297 26598
rect 14331 26564 14381 26598
rect 14247 26530 14381 26564
rect 14247 26496 14297 26530
rect 14331 26496 14381 26530
rect 14247 26462 14381 26496
rect 14247 26428 14297 26462
rect 14331 26428 14381 26462
rect 14247 26394 14381 26428
rect 14247 26360 14297 26394
rect 14331 26360 14381 26394
rect 14247 26326 14381 26360
rect 14247 26292 14297 26326
rect 14331 26292 14381 26326
rect 14247 26258 14381 26292
rect 14247 26224 14297 26258
rect 14331 26224 14381 26258
rect 14247 26190 14381 26224
rect 14247 26156 14297 26190
rect 14331 26156 14381 26190
rect 14247 26122 14381 26156
rect 14247 26088 14297 26122
rect 14331 26088 14381 26122
rect 14247 26054 14381 26088
rect 14247 26020 14297 26054
rect 14331 26020 14381 26054
rect 14247 25986 14381 26020
rect 14247 25952 14297 25986
rect 14331 25952 14381 25986
rect 14247 25918 14381 25952
rect 14247 25884 14297 25918
rect 14331 25884 14381 25918
rect 14247 25850 14381 25884
rect 14247 25816 14297 25850
rect 14331 25816 14381 25850
rect 14247 25782 14381 25816
rect 14247 25748 14297 25782
rect 14331 25748 14381 25782
rect 14247 25714 14381 25748
rect 14247 25680 14297 25714
rect 14331 25680 14381 25714
rect 14247 25646 14381 25680
rect 14247 25612 14297 25646
rect 14331 25612 14381 25646
rect 14247 25578 14381 25612
rect 14247 25544 14297 25578
rect 14331 25544 14381 25578
rect 14247 25510 14381 25544
rect 14247 25476 14297 25510
rect 14331 25476 14381 25510
rect 14247 25442 14381 25476
rect 14247 25408 14297 25442
rect 14331 25408 14381 25442
rect 14247 25374 14381 25408
rect 14247 25340 14297 25374
rect 14331 25340 14381 25374
rect 14247 25306 14381 25340
rect 14247 25272 14297 25306
rect 14331 25272 14381 25306
rect 14247 25238 14381 25272
rect 14247 25204 14297 25238
rect 14331 25204 14381 25238
rect 14247 25170 14381 25204
rect 14247 25136 14297 25170
rect 14331 25136 14381 25170
rect 14247 25102 14381 25136
rect 14247 25068 14297 25102
rect 14331 25068 14381 25102
rect 14247 25034 14381 25068
rect 14247 25000 14297 25034
rect 14331 25000 14381 25034
rect 14247 24966 14381 25000
rect 14247 24932 14297 24966
rect 14331 24932 14381 24966
rect 14247 24898 14381 24932
rect 14247 24864 14297 24898
rect 14331 24864 14381 24898
rect 14247 24830 14381 24864
rect 14247 24796 14297 24830
rect 14331 24796 14381 24830
rect 14247 24762 14381 24796
rect 14247 24728 14297 24762
rect 14331 24728 14381 24762
rect 14247 24694 14381 24728
rect 14247 24660 14297 24694
rect 14331 24660 14381 24694
rect 14247 24626 14381 24660
rect 14247 24592 14297 24626
rect 14331 24592 14381 24626
rect 14247 24558 14381 24592
rect 14247 24524 14297 24558
rect 14331 24524 14381 24558
rect 14247 24490 14381 24524
rect 14247 24456 14297 24490
rect 14331 24456 14381 24490
rect 14247 24422 14381 24456
rect 14247 24388 14297 24422
rect 14331 24388 14381 24422
rect 14247 24354 14381 24388
rect 14247 24320 14297 24354
rect 14331 24320 14381 24354
rect 14247 24286 14381 24320
rect 14247 24252 14297 24286
rect 14331 24252 14381 24286
rect 14247 24218 14381 24252
rect 14247 24184 14297 24218
rect 14331 24184 14381 24218
rect 14247 24150 14381 24184
rect 14247 24116 14297 24150
rect 14331 24116 14381 24150
rect 14247 24082 14381 24116
rect 14247 24048 14297 24082
rect 14331 24048 14381 24082
rect 14247 24014 14381 24048
rect 14247 23980 14297 24014
rect 14331 23980 14381 24014
rect 14247 23946 14381 23980
rect 14247 23912 14297 23946
rect 14331 23912 14381 23946
rect 14247 23878 14381 23912
rect 14247 23844 14297 23878
rect 14331 23844 14381 23878
rect 14247 23810 14381 23844
rect 14247 23776 14297 23810
rect 14331 23776 14381 23810
rect 14247 23742 14381 23776
rect 14247 23708 14297 23742
rect 14331 23708 14381 23742
rect 14247 23674 14381 23708
rect 14247 23640 14297 23674
rect 14331 23640 14381 23674
rect 14247 23606 14381 23640
rect 14247 23572 14297 23606
rect 14331 23572 14381 23606
rect 14247 23538 14381 23572
rect 14247 23504 14297 23538
rect 14331 23504 14381 23538
rect 14247 23470 14381 23504
rect 14247 23436 14297 23470
rect 14331 23436 14381 23470
rect 14247 23402 14381 23436
rect 14247 23368 14297 23402
rect 14331 23368 14381 23402
rect 14247 23334 14381 23368
rect 14247 23300 14297 23334
rect 14331 23300 14381 23334
rect 14247 23266 14381 23300
rect 14247 23232 14297 23266
rect 14331 23232 14381 23266
rect 14247 23198 14381 23232
rect 14247 23164 14297 23198
rect 14331 23164 14381 23198
rect 14247 23130 14381 23164
rect 14247 23096 14297 23130
rect 14331 23096 14381 23130
rect 14247 23062 14381 23096
rect 14247 23028 14297 23062
rect 14331 23028 14381 23062
rect 14247 22994 14381 23028
rect 14247 22960 14297 22994
rect 14331 22960 14381 22994
rect 14247 22926 14381 22960
rect 14247 22892 14297 22926
rect 14331 22892 14381 22926
rect 14247 22858 14381 22892
rect 14247 22824 14297 22858
rect 14331 22824 14381 22858
rect 14247 22790 14381 22824
rect 14247 22756 14297 22790
rect 14331 22756 14381 22790
rect 14247 22722 14381 22756
rect 14247 22688 14297 22722
rect 14331 22688 14381 22722
rect 14247 22654 14381 22688
rect 14247 22620 14297 22654
rect 14331 22620 14381 22654
rect 14247 22586 14381 22620
rect 14247 22552 14297 22586
rect 14331 22552 14381 22586
rect 14247 22518 14381 22552
rect 14247 22484 14297 22518
rect 14331 22484 14381 22518
rect 14247 22450 14381 22484
rect 14247 22416 14297 22450
rect 14331 22416 14381 22450
rect 14247 22382 14381 22416
rect 14247 22348 14297 22382
rect 14331 22348 14381 22382
rect 14247 22314 14381 22348
rect 14247 22280 14297 22314
rect 14331 22280 14381 22314
rect 14247 22246 14381 22280
rect 14247 22212 14297 22246
rect 14331 22212 14381 22246
rect 14247 22178 14381 22212
rect 14247 22144 14297 22178
rect 14331 22144 14381 22178
rect 14247 22110 14381 22144
rect 14247 22076 14297 22110
rect 14331 22076 14381 22110
rect 14247 22042 14381 22076
rect 14247 22008 14297 22042
rect 14331 22008 14381 22042
rect 14247 21974 14381 22008
rect 14247 21940 14297 21974
rect 14331 21940 14381 21974
rect 14247 21906 14381 21940
rect 14247 21872 14297 21906
rect 14331 21872 14381 21906
rect 14247 21838 14381 21872
rect 14247 21804 14297 21838
rect 14331 21804 14381 21838
rect 14247 21770 14381 21804
rect 14247 21736 14297 21770
rect 14331 21736 14381 21770
rect 14247 21702 14381 21736
rect 14247 21668 14297 21702
rect 14331 21668 14381 21702
rect 14247 21634 14381 21668
rect 14247 21600 14297 21634
rect 14331 21600 14381 21634
rect 14247 21566 14381 21600
rect 14247 21532 14297 21566
rect 14331 21532 14381 21566
rect 14247 21498 14381 21532
rect 14247 21464 14297 21498
rect 14331 21464 14381 21498
rect 14247 21430 14381 21464
rect 14247 21396 14297 21430
rect 14331 21396 14381 21430
rect 14247 21362 14381 21396
rect 14247 21328 14297 21362
rect 14331 21328 14381 21362
rect 14247 21294 14381 21328
rect 14247 21260 14297 21294
rect 14331 21260 14381 21294
rect 14247 21226 14381 21260
rect 14247 21192 14297 21226
rect 14331 21192 14381 21226
rect 14247 21158 14381 21192
rect 14247 21124 14297 21158
rect 14331 21124 14381 21158
rect 14247 21090 14381 21124
rect 14247 21056 14297 21090
rect 14331 21056 14381 21090
rect 14247 21022 14381 21056
rect 14247 20988 14297 21022
rect 14331 20988 14381 21022
rect 14247 20954 14381 20988
rect 14247 20920 14297 20954
rect 14331 20920 14381 20954
rect 14247 20886 14381 20920
rect 14247 20852 14297 20886
rect 14331 20852 14381 20886
rect 14247 20818 14381 20852
rect 14247 20784 14297 20818
rect 14331 20784 14381 20818
rect 14247 20750 14381 20784
rect 14247 20716 14297 20750
rect 14331 20716 14381 20750
rect 14247 20682 14381 20716
rect 14247 20648 14297 20682
rect 14331 20648 14381 20682
rect 14247 20614 14381 20648
rect 14247 20580 14297 20614
rect 14331 20580 14381 20614
rect 14247 20546 14381 20580
rect 14247 20512 14297 20546
rect 14331 20512 14381 20546
rect 14247 20478 14381 20512
rect 14247 20444 14297 20478
rect 14331 20444 14381 20478
rect 14247 20410 14381 20444
rect 14247 20376 14297 20410
rect 14331 20376 14381 20410
rect 14247 20342 14381 20376
rect 14247 20308 14297 20342
rect 14331 20308 14381 20342
rect 14247 20274 14381 20308
rect 14247 20240 14297 20274
rect 14331 20240 14381 20274
rect 14247 20206 14381 20240
rect 14247 20172 14297 20206
rect 14331 20172 14381 20206
rect 14247 20138 14381 20172
rect 14247 20104 14297 20138
rect 14331 20104 14381 20138
rect 14247 20070 14381 20104
rect 14247 20036 14297 20070
rect 14331 20036 14381 20070
rect 14247 20002 14381 20036
rect 14247 19968 14297 20002
rect 14331 19968 14381 20002
rect 14247 19934 14381 19968
rect 14247 19900 14297 19934
rect 14331 19900 14381 19934
rect 14247 19866 14381 19900
rect 14247 19832 14297 19866
rect 14331 19832 14381 19866
rect 14247 19798 14381 19832
rect 14247 19764 14297 19798
rect 14331 19764 14381 19798
rect 14247 19730 14381 19764
rect 14247 19696 14297 19730
rect 14331 19696 14381 19730
rect 14247 19662 14381 19696
rect 14247 19628 14297 19662
rect 14331 19628 14381 19662
rect 14247 19594 14381 19628
rect 14247 19560 14297 19594
rect 14331 19560 14381 19594
rect 14247 19526 14381 19560
rect 14247 19492 14297 19526
rect 14331 19492 14381 19526
rect 14247 19458 14381 19492
rect 14247 19424 14297 19458
rect 14331 19424 14381 19458
rect 14247 19390 14381 19424
rect 14247 19356 14297 19390
rect 14331 19356 14381 19390
rect 14247 19322 14381 19356
rect 14247 19288 14297 19322
rect 14331 19288 14381 19322
rect 14247 19254 14381 19288
rect 14247 19220 14297 19254
rect 14331 19220 14381 19254
rect 14247 19186 14381 19220
rect 14247 19152 14297 19186
rect 14331 19152 14381 19186
rect 14247 19118 14381 19152
rect 14247 19084 14297 19118
rect 14331 19084 14381 19118
rect 14247 19050 14381 19084
rect 14247 19016 14297 19050
rect 14331 19016 14381 19050
rect 14247 18982 14381 19016
rect 14247 18948 14297 18982
rect 14331 18948 14381 18982
rect 14247 18914 14381 18948
rect 14247 18880 14297 18914
rect 14331 18880 14381 18914
rect 14247 18846 14381 18880
rect 14247 18812 14297 18846
rect 14331 18812 14381 18846
rect 14247 18778 14381 18812
rect 14247 18744 14297 18778
rect 14331 18744 14381 18778
rect 14247 18710 14381 18744
rect 14247 18676 14297 18710
rect 14331 18676 14381 18710
rect 14247 18642 14381 18676
rect 14247 18608 14297 18642
rect 14331 18608 14381 18642
rect 14247 18574 14381 18608
rect 14247 18540 14297 18574
rect 14331 18540 14381 18574
rect 14247 18506 14381 18540
rect 14247 18472 14297 18506
rect 14331 18472 14381 18506
rect 14247 18438 14381 18472
rect 14247 18404 14297 18438
rect 14331 18404 14381 18438
rect 14247 18370 14381 18404
rect 14247 18336 14297 18370
rect 14331 18336 14381 18370
rect 14247 18302 14381 18336
rect 14247 18268 14297 18302
rect 14331 18268 14381 18302
rect 14247 18234 14381 18268
rect 14247 18200 14297 18234
rect 14331 18200 14381 18234
rect 14247 18166 14381 18200
rect 14247 18132 14297 18166
rect 14331 18132 14381 18166
rect 14247 18098 14381 18132
rect 14247 18064 14297 18098
rect 14331 18064 14381 18098
rect 14247 18030 14381 18064
rect 14247 17996 14297 18030
rect 14331 17996 14381 18030
rect 14247 17962 14381 17996
rect 14247 17928 14297 17962
rect 14331 17928 14381 17962
rect 14247 17894 14381 17928
rect 14247 17860 14297 17894
rect 14331 17860 14381 17894
rect 14247 17826 14381 17860
rect 14247 17792 14297 17826
rect 14331 17792 14381 17826
rect 14247 17758 14381 17792
rect 14247 17724 14297 17758
rect 14331 17724 14381 17758
rect 14247 17690 14381 17724
rect 14247 17656 14297 17690
rect 14331 17656 14381 17690
rect 14247 17622 14381 17656
rect 14247 17588 14297 17622
rect 14331 17588 14381 17622
rect 14247 17554 14381 17588
rect 14247 17520 14297 17554
rect 14331 17520 14381 17554
rect 14247 17486 14381 17520
rect 14247 17452 14297 17486
rect 14331 17452 14381 17486
rect 14247 17418 14381 17452
rect 14247 17384 14297 17418
rect 14331 17384 14381 17418
rect 14247 17350 14381 17384
rect 14247 17316 14297 17350
rect 14331 17316 14381 17350
rect 14247 17282 14381 17316
rect 14247 17248 14297 17282
rect 14331 17248 14381 17282
rect 14247 17214 14381 17248
rect 14247 17180 14297 17214
rect 14331 17180 14381 17214
rect 14247 17146 14381 17180
rect 14247 17112 14297 17146
rect 14331 17112 14381 17146
rect 14247 17078 14381 17112
rect 14247 17044 14297 17078
rect 14331 17044 14381 17078
rect 14247 17010 14381 17044
rect 14247 16976 14297 17010
rect 14331 16976 14381 17010
rect 14247 16942 14381 16976
rect 14247 16908 14297 16942
rect 14331 16908 14381 16942
rect 14247 16874 14381 16908
rect 14247 16840 14297 16874
rect 14331 16840 14381 16874
rect 14247 16806 14381 16840
rect 14247 16772 14297 16806
rect 14331 16772 14381 16806
rect 14247 16738 14381 16772
rect 14247 16704 14297 16738
rect 14331 16704 14381 16738
rect 14247 16670 14381 16704
rect 14247 16636 14297 16670
rect 14331 16636 14381 16670
rect 14247 16602 14381 16636
rect 14247 16568 14297 16602
rect 14331 16568 14381 16602
rect 14247 16534 14381 16568
rect 14247 16500 14297 16534
rect 14331 16500 14381 16534
rect 14247 16466 14381 16500
rect 14247 16432 14297 16466
rect 14331 16432 14381 16466
rect 14247 16398 14381 16432
rect 14247 16364 14297 16398
rect 14331 16364 14381 16398
rect 14247 16330 14381 16364
rect 14247 16296 14297 16330
rect 14331 16296 14381 16330
rect 14247 16262 14381 16296
rect 14247 16228 14297 16262
rect 14331 16228 14381 16262
rect 14247 16194 14381 16228
rect 14247 16160 14297 16194
rect 14331 16160 14381 16194
rect 14247 16126 14381 16160
rect 14247 16092 14297 16126
rect 14331 16092 14381 16126
rect 14247 16058 14381 16092
rect 14247 16024 14297 16058
rect 14331 16024 14381 16058
rect 14247 15990 14381 16024
rect 14247 15956 14297 15990
rect 14331 15956 14381 15990
rect 14247 15922 14381 15956
rect 14247 15888 14297 15922
rect 14331 15888 14381 15922
rect 14247 15854 14381 15888
rect 14247 15820 14297 15854
rect 14331 15820 14381 15854
rect 14247 15786 14381 15820
rect 14247 15752 14297 15786
rect 14331 15752 14381 15786
rect 14247 15718 14381 15752
rect 14247 15684 14297 15718
rect 14331 15684 14381 15718
rect 14247 15650 14381 15684
rect 14247 15616 14297 15650
rect 14331 15616 14381 15650
rect 14247 15582 14381 15616
rect 14247 15548 14297 15582
rect 14331 15548 14381 15582
rect 14247 15514 14381 15548
rect 14247 15480 14297 15514
rect 14331 15480 14381 15514
rect 14247 15446 14381 15480
rect 14247 15412 14297 15446
rect 14331 15412 14381 15446
rect 14247 15378 14381 15412
rect 14247 15344 14297 15378
rect 14331 15344 14381 15378
rect 14247 15310 14381 15344
rect 14247 15276 14297 15310
rect 14331 15276 14381 15310
rect 14247 15242 14381 15276
rect 14247 15208 14297 15242
rect 14331 15208 14381 15242
rect 583 15140 632 15174
rect 666 15140 715 15174
rect 583 15106 715 15140
rect 583 15072 632 15106
rect 666 15072 715 15106
rect 583 15038 715 15072
rect 583 15004 632 15038
rect 666 15004 715 15038
rect 583 14970 715 15004
rect 583 14936 632 14970
rect 666 14936 715 14970
rect 583 14902 715 14936
rect 583 14868 632 14902
rect 666 14868 715 14902
rect 583 14825 715 14868
rect 14247 15174 14381 15208
rect 14247 15140 14297 15174
rect 14331 15140 14381 15174
rect 14247 15106 14381 15140
rect 14247 15072 14297 15106
rect 14331 15072 14381 15106
rect 14247 15038 14381 15072
rect 14247 15004 14297 15038
rect 14331 15004 14381 15038
rect 14247 14970 14381 15004
rect 14247 14936 14297 14970
rect 14331 14936 14381 14970
rect 14247 14902 14381 14936
rect 14247 14868 14297 14902
rect 14331 14868 14381 14902
rect 14247 14825 14381 14868
rect 583 14775 14381 14825
rect 583 14741 766 14775
rect 800 14741 834 14775
rect 868 14741 902 14775
rect 936 14741 970 14775
rect 1004 14741 1038 14775
rect 1072 14741 1106 14775
rect 1140 14741 1174 14775
rect 1208 14741 1242 14775
rect 1276 14741 1310 14775
rect 1344 14741 1378 14775
rect 1412 14741 1446 14775
rect 1480 14741 1514 14775
rect 1548 14741 1582 14775
rect 1616 14741 1650 14775
rect 1684 14741 1718 14775
rect 1752 14741 1786 14775
rect 1820 14741 1854 14775
rect 1888 14741 1922 14775
rect 1956 14741 1990 14775
rect 2024 14741 2058 14775
rect 2092 14741 2126 14775
rect 2160 14741 2194 14775
rect 2228 14741 2262 14775
rect 2296 14741 2330 14775
rect 2364 14741 2398 14775
rect 2432 14741 2466 14775
rect 2500 14741 2534 14775
rect 2568 14741 2602 14775
rect 2636 14741 2670 14775
rect 2704 14741 2738 14775
rect 2772 14741 2806 14775
rect 2840 14741 2874 14775
rect 2908 14741 2942 14775
rect 2976 14741 3010 14775
rect 3044 14741 3078 14775
rect 3112 14741 3146 14775
rect 3180 14741 3214 14775
rect 3248 14741 3282 14775
rect 3316 14741 3350 14775
rect 3384 14741 3418 14775
rect 3452 14741 3486 14775
rect 3520 14741 3554 14775
rect 3588 14741 3622 14775
rect 3656 14741 3690 14775
rect 3724 14741 3758 14775
rect 3792 14741 3826 14775
rect 3860 14741 3894 14775
rect 3928 14741 3962 14775
rect 3996 14741 4030 14775
rect 4064 14741 4098 14775
rect 4132 14741 4166 14775
rect 4200 14741 4234 14775
rect 4268 14741 4302 14775
rect 4336 14741 4370 14775
rect 4404 14741 4438 14775
rect 4472 14741 4506 14775
rect 4540 14741 4574 14775
rect 4608 14741 4642 14775
rect 4676 14741 4710 14775
rect 4744 14741 4778 14775
rect 4812 14741 4846 14775
rect 4880 14741 4914 14775
rect 4948 14741 4982 14775
rect 5016 14741 5050 14775
rect 5084 14741 5118 14775
rect 5152 14741 5186 14775
rect 5220 14741 5254 14775
rect 5288 14741 5322 14775
rect 5356 14741 5390 14775
rect 5424 14741 5458 14775
rect 5492 14741 5526 14775
rect 5560 14741 5594 14775
rect 5628 14741 5662 14775
rect 5696 14741 5730 14775
rect 5764 14741 5798 14775
rect 5832 14741 5866 14775
rect 5900 14741 5934 14775
rect 5968 14741 6002 14775
rect 6036 14741 6070 14775
rect 6104 14741 6138 14775
rect 6172 14741 6206 14775
rect 6240 14741 6274 14775
rect 6308 14741 6342 14775
rect 6376 14741 6410 14775
rect 6444 14741 6478 14775
rect 6512 14741 6546 14775
rect 6580 14741 6614 14775
rect 6648 14741 6682 14775
rect 6716 14741 6750 14775
rect 6784 14741 6818 14775
rect 6852 14741 6886 14775
rect 6920 14741 6954 14775
rect 6988 14741 7022 14775
rect 7056 14741 7090 14775
rect 7124 14741 7158 14775
rect 7192 14741 7226 14775
rect 7260 14741 7294 14775
rect 7328 14741 7362 14775
rect 7396 14741 7430 14775
rect 7464 14741 7498 14775
rect 7532 14741 7566 14775
rect 7600 14741 7634 14775
rect 7668 14741 7702 14775
rect 7736 14741 7770 14775
rect 7804 14741 7838 14775
rect 7872 14741 7906 14775
rect 7940 14741 7974 14775
rect 8008 14741 8042 14775
rect 8076 14741 8110 14775
rect 8144 14741 8178 14775
rect 8212 14741 8246 14775
rect 8280 14741 8314 14775
rect 8348 14741 8382 14775
rect 8416 14741 8450 14775
rect 8484 14741 8518 14775
rect 8552 14741 8586 14775
rect 8620 14741 8654 14775
rect 8688 14741 8722 14775
rect 8756 14741 8790 14775
rect 8824 14741 8858 14775
rect 8892 14741 8926 14775
rect 8960 14741 8994 14775
rect 9028 14741 9062 14775
rect 9096 14741 9130 14775
rect 9164 14741 9198 14775
rect 9232 14741 9266 14775
rect 9300 14741 9334 14775
rect 9368 14741 9402 14775
rect 9436 14741 9470 14775
rect 9504 14741 9538 14775
rect 9572 14741 9606 14775
rect 9640 14741 9674 14775
rect 9708 14741 9742 14775
rect 9776 14741 9810 14775
rect 9844 14741 9878 14775
rect 9912 14741 9946 14775
rect 9980 14741 10014 14775
rect 10048 14741 10082 14775
rect 10116 14741 10150 14775
rect 10184 14741 10218 14775
rect 10252 14741 10286 14775
rect 10320 14741 10354 14775
rect 10388 14741 10422 14775
rect 10456 14741 10490 14775
rect 10524 14741 10558 14775
rect 10592 14741 10626 14775
rect 10660 14741 10694 14775
rect 10728 14741 10762 14775
rect 10796 14741 10830 14775
rect 10864 14741 10898 14775
rect 10932 14741 10966 14775
rect 11000 14741 11034 14775
rect 11068 14741 11102 14775
rect 11136 14741 11170 14775
rect 11204 14741 11238 14775
rect 11272 14741 11306 14775
rect 11340 14741 11374 14775
rect 11408 14741 11442 14775
rect 11476 14741 11510 14775
rect 11544 14741 11578 14775
rect 11612 14741 11646 14775
rect 11680 14741 11714 14775
rect 11748 14741 11782 14775
rect 11816 14741 11850 14775
rect 11884 14741 11918 14775
rect 11952 14741 11986 14775
rect 12020 14741 12054 14775
rect 12088 14741 12122 14775
rect 12156 14741 12190 14775
rect 12224 14741 12258 14775
rect 12292 14741 12326 14775
rect 12360 14741 12394 14775
rect 12428 14741 12462 14775
rect 12496 14741 12530 14775
rect 12564 14741 12598 14775
rect 12632 14741 12666 14775
rect 12700 14741 12734 14775
rect 12768 14741 12802 14775
rect 12836 14741 12870 14775
rect 12904 14741 12938 14775
rect 12972 14741 13006 14775
rect 13040 14741 13074 14775
rect 13108 14741 13142 14775
rect 13176 14741 13210 14775
rect 13244 14741 13278 14775
rect 13312 14741 13346 14775
rect 13380 14741 13414 14775
rect 13448 14741 13482 14775
rect 13516 14741 13550 14775
rect 13584 14741 13618 14775
rect 13652 14741 13686 14775
rect 13720 14741 13754 14775
rect 13788 14741 13822 14775
rect 13856 14741 13890 14775
rect 13924 14741 13958 14775
rect 13992 14741 14026 14775
rect 14060 14741 14094 14775
rect 14128 14741 14162 14775
rect 14196 14741 14381 14775
rect 583 14691 14381 14741
<< mvpsubdiffcont >>
rect 455 36463 489 36497
rect 523 36463 557 36497
rect 591 36463 625 36497
rect 659 36463 693 36497
rect 727 36463 761 36497
rect 795 36463 829 36497
rect 863 36463 897 36497
rect 931 36463 965 36497
rect 999 36463 1033 36497
rect 1067 36463 1101 36497
rect 1135 36463 1169 36497
rect 1203 36463 1237 36497
rect 1271 36463 1305 36497
rect 1339 36463 1373 36497
rect 1407 36463 1441 36497
rect 1475 36463 1509 36497
rect 1543 36463 1577 36497
rect 1611 36463 1645 36497
rect 1679 36463 1713 36497
rect 1747 36463 1781 36497
rect 1815 36463 1849 36497
rect 1883 36463 1917 36497
rect 1951 36463 1985 36497
rect 2019 36463 2053 36497
rect 2087 36463 2121 36497
rect 2155 36463 2189 36497
rect 2223 36463 2257 36497
rect 2291 36463 2325 36497
rect 2359 36463 2393 36497
rect 2427 36463 2461 36497
rect 2495 36463 2529 36497
rect 2563 36463 2597 36497
rect 2631 36463 2665 36497
rect 2699 36463 2733 36497
rect 2767 36463 2801 36497
rect 2835 36463 2869 36497
rect 2903 36463 2937 36497
rect 2971 36463 3005 36497
rect 3039 36463 3073 36497
rect 3107 36463 3141 36497
rect 3175 36463 3209 36497
rect 3243 36463 3277 36497
rect 3311 36463 3345 36497
rect 3379 36463 3413 36497
rect 3447 36463 3481 36497
rect 3515 36463 3549 36497
rect 3583 36463 3617 36497
rect 3651 36463 3685 36497
rect 3719 36463 3753 36497
rect 3787 36463 3821 36497
rect 3855 36463 3889 36497
rect 3923 36463 3957 36497
rect 3991 36463 4025 36497
rect 4059 36463 4093 36497
rect 4127 36463 4161 36497
rect 4195 36463 4229 36497
rect 4263 36463 4297 36497
rect 4331 36463 4365 36497
rect 4399 36463 4433 36497
rect 4467 36463 4501 36497
rect 4535 36463 4569 36497
rect 4603 36463 4637 36497
rect 4671 36463 4705 36497
rect 4739 36463 4773 36497
rect 4807 36463 4841 36497
rect 4875 36463 4909 36497
rect 4943 36463 4977 36497
rect 5011 36463 5045 36497
rect 5079 36463 5113 36497
rect 5147 36463 5181 36497
rect 5215 36463 5249 36497
rect 5283 36463 5317 36497
rect 5351 36463 5385 36497
rect 5419 36463 5453 36497
rect 5487 36463 5521 36497
rect 5555 36463 5589 36497
rect 5623 36463 5657 36497
rect 5691 36463 5725 36497
rect 5759 36463 5793 36497
rect 5827 36463 5861 36497
rect 5895 36463 5929 36497
rect 5963 36463 5997 36497
rect 6031 36463 6065 36497
rect 6099 36463 6133 36497
rect 6167 36463 6201 36497
rect 6235 36463 6269 36497
rect 6303 36463 6337 36497
rect 6371 36463 6405 36497
rect 6439 36463 6473 36497
rect 6507 36463 6541 36497
rect 6575 36463 6609 36497
rect 6643 36463 6677 36497
rect 6711 36463 6745 36497
rect 6779 36463 6813 36497
rect 6847 36463 6881 36497
rect 6915 36463 6949 36497
rect 6983 36463 7017 36497
rect 7051 36463 7085 36497
rect 7119 36463 7153 36497
rect 7187 36463 7221 36497
rect 7255 36463 7289 36497
rect 7323 36463 7357 36497
rect 7391 36463 7425 36497
rect 7459 36463 7493 36497
rect 7527 36463 7561 36497
rect 7595 36463 7629 36497
rect 7663 36463 7697 36497
rect 7731 36463 7765 36497
rect 7799 36463 7833 36497
rect 7867 36463 7901 36497
rect 7935 36463 7969 36497
rect 8003 36463 8037 36497
rect 8071 36463 8105 36497
rect 8139 36463 8173 36497
rect 8207 36463 8241 36497
rect 8275 36463 8309 36497
rect 8343 36463 8377 36497
rect 8411 36463 8445 36497
rect 8479 36463 8513 36497
rect 8547 36463 8581 36497
rect 8615 36463 8649 36497
rect 8683 36463 8717 36497
rect 8751 36463 8785 36497
rect 8819 36463 8853 36497
rect 8887 36463 8921 36497
rect 8955 36463 8989 36497
rect 9023 36463 9057 36497
rect 9091 36463 9125 36497
rect 9159 36463 9193 36497
rect 9227 36463 9261 36497
rect 9295 36463 9329 36497
rect 9363 36463 9397 36497
rect 9431 36463 9465 36497
rect 9499 36463 9533 36497
rect 9567 36463 9601 36497
rect 9635 36463 9669 36497
rect 9703 36463 9737 36497
rect 9771 36463 9805 36497
rect 9839 36463 9873 36497
rect 9907 36463 9941 36497
rect 9975 36463 10009 36497
rect 10043 36463 10077 36497
rect 10111 36463 10145 36497
rect 10179 36463 10213 36497
rect 10247 36463 10281 36497
rect 10315 36463 10349 36497
rect 10383 36463 10417 36497
rect 10451 36463 10485 36497
rect 10519 36463 10553 36497
rect 10587 36463 10621 36497
rect 10655 36463 10689 36497
rect 10723 36463 10757 36497
rect 10791 36463 10825 36497
rect 10859 36463 10893 36497
rect 10927 36463 10961 36497
rect 10995 36463 11029 36497
rect 11063 36463 11097 36497
rect 11131 36463 11165 36497
rect 11199 36463 11233 36497
rect 11267 36463 11301 36497
rect 11335 36463 11369 36497
rect 11403 36463 11437 36497
rect 11471 36463 11505 36497
rect 11539 36463 11573 36497
rect 11607 36463 11641 36497
rect 11675 36463 11709 36497
rect 11743 36463 11777 36497
rect 11811 36463 11845 36497
rect 11879 36463 11913 36497
rect 11947 36463 11981 36497
rect 12015 36463 12049 36497
rect 12083 36463 12117 36497
rect 12151 36463 12185 36497
rect 12219 36463 12253 36497
rect 12287 36463 12321 36497
rect 12355 36463 12389 36497
rect 12423 36463 12457 36497
rect 12491 36463 12525 36497
rect 12559 36463 12593 36497
rect 12627 36463 12661 36497
rect 12695 36463 12729 36497
rect 12763 36463 12797 36497
rect 12831 36463 12865 36497
rect 12899 36463 12933 36497
rect 12967 36463 13001 36497
rect 13035 36463 13069 36497
rect 13103 36463 13137 36497
rect 13171 36463 13205 36497
rect 13239 36463 13273 36497
rect 13307 36463 13341 36497
rect 13375 36463 13409 36497
rect 13443 36463 13477 36497
rect 13511 36463 13545 36497
rect 13579 36463 13613 36497
rect 13647 36463 13681 36497
rect 13715 36463 13749 36497
rect 13783 36463 13817 36497
rect 13851 36463 13885 36497
rect 13919 36463 13953 36497
rect 13987 36463 14021 36497
rect 14055 36463 14089 36497
rect 14123 36463 14157 36497
rect 14191 36463 14225 36497
rect 14259 36463 14293 36497
rect 14327 36463 14361 36497
rect 14395 36463 14429 36497
rect 14463 36463 14497 36497
rect 312 36322 346 36356
rect 312 36254 346 36288
rect 14607 36328 14641 36362
rect 14607 36260 14641 36294
rect 312 36186 346 36220
rect 312 36118 346 36152
rect 312 36050 346 36084
rect 312 35982 346 36016
rect 312 35914 346 35948
rect 312 35846 346 35880
rect 312 35778 346 35812
rect 312 35710 346 35744
rect 312 35642 346 35676
rect 312 35574 346 35608
rect 312 35506 346 35540
rect 312 35438 346 35472
rect 312 35370 346 35404
rect 312 35302 346 35336
rect 312 35234 346 35268
rect 312 35166 346 35200
rect 312 35098 346 35132
rect 312 35030 346 35064
rect 312 34962 346 34996
rect 312 34894 346 34928
rect 312 34826 346 34860
rect 312 34758 346 34792
rect 312 34690 346 34724
rect 312 34622 346 34656
rect 312 34554 346 34588
rect 312 34486 346 34520
rect 312 34418 346 34452
rect 312 34350 346 34384
rect 312 34282 346 34316
rect 312 34214 346 34248
rect 312 34146 346 34180
rect 312 34078 346 34112
rect 312 34010 346 34044
rect 312 33942 346 33976
rect 312 33874 346 33908
rect 312 33806 346 33840
rect 312 33738 346 33772
rect 312 33670 346 33704
rect 312 33602 346 33636
rect 312 33534 346 33568
rect 312 33466 346 33500
rect 312 33398 346 33432
rect 312 33330 346 33364
rect 312 33262 346 33296
rect 312 33194 346 33228
rect 312 33126 346 33160
rect 312 33058 346 33092
rect 312 32990 346 33024
rect 312 32922 346 32956
rect 312 32854 346 32888
rect 312 32786 346 32820
rect 312 32718 346 32752
rect 312 32650 346 32684
rect 312 32582 346 32616
rect 312 32514 346 32548
rect 312 32446 346 32480
rect 312 32378 346 32412
rect 312 32310 346 32344
rect 312 32242 346 32276
rect 312 32174 346 32208
rect 312 32106 346 32140
rect 312 32038 346 32072
rect 312 31970 346 32004
rect 312 31902 346 31936
rect 312 31834 346 31868
rect 312 31766 346 31800
rect 312 31698 346 31732
rect 312 31630 346 31664
rect 312 31562 346 31596
rect 312 31494 346 31528
rect 312 31426 346 31460
rect 312 31358 346 31392
rect 312 31290 346 31324
rect 312 31222 346 31256
rect 312 31154 346 31188
rect 312 31086 346 31120
rect 312 31018 346 31052
rect 312 30950 346 30984
rect 312 30882 346 30916
rect 312 30814 346 30848
rect 312 30746 346 30780
rect 312 30678 346 30712
rect 312 30610 346 30644
rect 312 30542 346 30576
rect 312 30474 346 30508
rect 312 30406 346 30440
rect 312 30338 346 30372
rect 312 30270 346 30304
rect 312 30202 346 30236
rect 312 30134 346 30168
rect 312 30066 346 30100
rect 312 29998 346 30032
rect 312 29930 346 29964
rect 312 29862 346 29896
rect 312 29794 346 29828
rect 312 29726 346 29760
rect 312 29658 346 29692
rect 312 29590 346 29624
rect 312 29522 346 29556
rect 312 29454 346 29488
rect 312 29386 346 29420
rect 312 29318 346 29352
rect 312 29250 346 29284
rect 312 29182 346 29216
rect 312 29114 346 29148
rect 312 29046 346 29080
rect 312 28978 346 29012
rect 312 28910 346 28944
rect 312 28842 346 28876
rect 312 28774 346 28808
rect 312 28706 346 28740
rect 312 28638 346 28672
rect 312 28570 346 28604
rect 312 28502 346 28536
rect 312 28434 346 28468
rect 312 28366 346 28400
rect 312 28298 346 28332
rect 312 28230 346 28264
rect 312 28162 346 28196
rect 312 28094 346 28128
rect 312 28026 346 28060
rect 312 27958 346 27992
rect 312 27890 346 27924
rect 312 27822 346 27856
rect 312 27754 346 27788
rect 312 27686 346 27720
rect 312 27618 346 27652
rect 312 27550 346 27584
rect 312 27482 346 27516
rect 312 27414 346 27448
rect 312 27346 346 27380
rect 312 27278 346 27312
rect 312 27210 346 27244
rect 312 27142 346 27176
rect 312 27074 346 27108
rect 312 27006 346 27040
rect 312 26938 346 26972
rect 312 26870 346 26904
rect 312 26802 346 26836
rect 312 26734 346 26768
rect 312 26666 346 26700
rect 312 26598 346 26632
rect 312 26530 346 26564
rect 312 26462 346 26496
rect 312 26394 346 26428
rect 312 26326 346 26360
rect 312 26258 346 26292
rect 312 26190 346 26224
rect 312 26122 346 26156
rect 312 26054 346 26088
rect 312 25986 346 26020
rect 312 25918 346 25952
rect 312 25850 346 25884
rect 312 25782 346 25816
rect 312 25714 346 25748
rect 312 25646 346 25680
rect 312 25578 346 25612
rect 312 25510 346 25544
rect 312 25442 346 25476
rect 312 25374 346 25408
rect 312 25306 346 25340
rect 312 25238 346 25272
rect 312 25170 346 25204
rect 312 25102 346 25136
rect 312 25034 346 25068
rect 312 24966 346 25000
rect 312 24898 346 24932
rect 312 24830 346 24864
rect 312 24762 346 24796
rect 312 24694 346 24728
rect 312 24626 346 24660
rect 312 24558 346 24592
rect 312 24490 346 24524
rect 312 24422 346 24456
rect 312 24354 346 24388
rect 312 24286 346 24320
rect 312 24218 346 24252
rect 312 24150 346 24184
rect 312 24082 346 24116
rect 312 24014 346 24048
rect 312 23946 346 23980
rect 312 23878 346 23912
rect 312 23810 346 23844
rect 312 23742 346 23776
rect 312 23674 346 23708
rect 312 23606 346 23640
rect 312 23538 346 23572
rect 312 23470 346 23504
rect 312 23402 346 23436
rect 312 23334 346 23368
rect 312 23266 346 23300
rect 312 23198 346 23232
rect 312 23130 346 23164
rect 312 23062 346 23096
rect 312 22994 346 23028
rect 312 22926 346 22960
rect 312 22858 346 22892
rect 312 22790 346 22824
rect 312 22722 346 22756
rect 312 22654 346 22688
rect 312 22586 346 22620
rect 312 22518 346 22552
rect 312 22450 346 22484
rect 312 22382 346 22416
rect 312 22314 346 22348
rect 312 22246 346 22280
rect 312 22178 346 22212
rect 312 22110 346 22144
rect 312 22042 346 22076
rect 312 21974 346 22008
rect 312 21906 346 21940
rect 312 21838 346 21872
rect 312 21770 346 21804
rect 312 21702 346 21736
rect 312 21634 346 21668
rect 312 21566 346 21600
rect 312 21498 346 21532
rect 312 21430 346 21464
rect 312 21362 346 21396
rect 312 21294 346 21328
rect 312 21226 346 21260
rect 312 21158 346 21192
rect 312 21090 346 21124
rect 312 21022 346 21056
rect 312 20954 346 20988
rect 312 20886 346 20920
rect 312 20818 346 20852
rect 312 20750 346 20784
rect 312 20682 346 20716
rect 312 20614 346 20648
rect 312 20546 346 20580
rect 312 20478 346 20512
rect 312 20410 346 20444
rect 312 20342 346 20376
rect 312 20274 346 20308
rect 312 20206 346 20240
rect 312 20138 346 20172
rect 312 20070 346 20104
rect 312 20002 346 20036
rect 312 19934 346 19968
rect 312 19866 346 19900
rect 312 19798 346 19832
rect 312 19730 346 19764
rect 312 19662 346 19696
rect 312 19594 346 19628
rect 312 19526 346 19560
rect 312 19458 346 19492
rect 312 19390 346 19424
rect 312 19322 346 19356
rect 312 19254 346 19288
rect 312 19186 346 19220
rect 312 19118 346 19152
rect 312 19050 346 19084
rect 312 18982 346 19016
rect 312 18914 346 18948
rect 312 18846 346 18880
rect 312 18778 346 18812
rect 312 18710 346 18744
rect 312 18642 346 18676
rect 312 18574 346 18608
rect 312 18506 346 18540
rect 312 18438 346 18472
rect 312 18370 346 18404
rect 312 18302 346 18336
rect 312 18234 346 18268
rect 312 18166 346 18200
rect 312 18098 346 18132
rect 312 18030 346 18064
rect 312 17962 346 17996
rect 312 17894 346 17928
rect 312 17826 346 17860
rect 312 17758 346 17792
rect 312 17690 346 17724
rect 312 17622 346 17656
rect 312 17554 346 17588
rect 312 17486 346 17520
rect 312 17418 346 17452
rect 312 17350 346 17384
rect 312 17282 346 17316
rect 312 17214 346 17248
rect 312 17146 346 17180
rect 312 17078 346 17112
rect 312 17010 346 17044
rect 312 16942 346 16976
rect 312 16874 346 16908
rect 312 16806 346 16840
rect 312 16738 346 16772
rect 312 16670 346 16704
rect 312 16602 346 16636
rect 312 16534 346 16568
rect 312 16466 346 16500
rect 312 16398 346 16432
rect 312 16330 346 16364
rect 312 16262 346 16296
rect 312 16194 346 16228
rect 312 16126 346 16160
rect 312 16058 346 16092
rect 312 15990 346 16024
rect 312 15922 346 15956
rect 312 15854 346 15888
rect 312 15786 346 15820
rect 312 15718 346 15752
rect 312 15650 346 15684
rect 312 15582 346 15616
rect 312 15514 346 15548
rect 312 15446 346 15480
rect 312 15378 346 15412
rect 312 15310 346 15344
rect 312 15242 346 15276
rect 312 15174 346 15208
rect 312 15106 346 15140
rect 312 15038 346 15072
rect 312 14970 346 15004
rect 312 14902 346 14936
rect 312 14834 346 14868
rect 312 14766 346 14800
rect 312 14698 346 14732
rect 1305 34645 1339 34679
rect 1373 34645 1407 34679
rect 1441 34645 1475 34679
rect 1509 34645 1543 34679
rect 1577 34645 1611 34679
rect 1645 34645 1679 34679
rect 1713 34645 1747 34679
rect 1781 34645 1815 34679
rect 1849 34645 1883 34679
rect 1917 34645 1951 34679
rect 1985 34645 2019 34679
rect 2053 34645 2087 34679
rect 2121 34645 2155 34679
rect 2189 34645 2223 34679
rect 2257 34645 2291 34679
rect 2325 34645 2359 34679
rect 2393 34645 2427 34679
rect 2461 34645 2495 34679
rect 2529 34645 2563 34679
rect 2597 34645 2631 34679
rect 2665 34645 2699 34679
rect 2733 34645 2767 34679
rect 2801 34645 2835 34679
rect 2869 34645 2903 34679
rect 2937 34645 2971 34679
rect 3005 34645 3039 34679
rect 3073 34645 3107 34679
rect 3141 34645 3175 34679
rect 3209 34645 3243 34679
rect 3277 34645 3311 34679
rect 3345 34645 3379 34679
rect 3413 34645 3447 34679
rect 3481 34645 3515 34679
rect 3549 34645 3583 34679
rect 3617 34645 3651 34679
rect 3685 34645 3719 34679
rect 3753 34645 3787 34679
rect 3821 34645 3855 34679
rect 3889 34645 3923 34679
rect 3957 34645 3991 34679
rect 4025 34645 4059 34679
rect 4093 34645 4127 34679
rect 4161 34645 4195 34679
rect 4229 34645 4263 34679
rect 4297 34645 4331 34679
rect 4365 34645 4399 34679
rect 4433 34645 4467 34679
rect 4501 34645 4535 34679
rect 4569 34645 4603 34679
rect 4637 34645 4671 34679
rect 4705 34645 4739 34679
rect 4773 34645 4807 34679
rect 4841 34645 4875 34679
rect 4909 34645 4943 34679
rect 4977 34645 5011 34679
rect 5045 34645 5079 34679
rect 5113 34645 5147 34679
rect 5181 34645 5215 34679
rect 5249 34645 5283 34679
rect 5317 34645 5351 34679
rect 5385 34645 5419 34679
rect 5453 34645 5487 34679
rect 5521 34645 5555 34679
rect 5589 34645 5623 34679
rect 5657 34645 5691 34679
rect 5725 34645 5759 34679
rect 5793 34645 5827 34679
rect 5861 34645 5895 34679
rect 5929 34645 5963 34679
rect 5997 34645 6031 34679
rect 6065 34645 6099 34679
rect 6133 34645 6167 34679
rect 6201 34645 6235 34679
rect 6269 34645 6303 34679
rect 6337 34645 6371 34679
rect 6405 34645 6439 34679
rect 6473 34645 6507 34679
rect 6541 34645 6575 34679
rect 6609 34645 6643 34679
rect 6677 34645 6711 34679
rect 6745 34645 6779 34679
rect 6813 34645 6847 34679
rect 6881 34645 6915 34679
rect 6949 34645 6983 34679
rect 7017 34645 7051 34679
rect 7085 34645 7119 34679
rect 7153 34645 7187 34679
rect 7221 34645 7255 34679
rect 7289 34645 7323 34679
rect 7357 34645 7391 34679
rect 7425 34645 7459 34679
rect 7493 34645 7527 34679
rect 7561 34645 7595 34679
rect 7629 34645 7663 34679
rect 7697 34645 7731 34679
rect 7765 34645 7799 34679
rect 7833 34645 7867 34679
rect 7901 34645 7935 34679
rect 7969 34645 8003 34679
rect 8037 34645 8071 34679
rect 8105 34645 8139 34679
rect 8173 34645 8207 34679
rect 8241 34645 8275 34679
rect 8309 34645 8343 34679
rect 8377 34645 8411 34679
rect 8445 34645 8479 34679
rect 8513 34645 8547 34679
rect 8581 34645 8615 34679
rect 8649 34645 8683 34679
rect 8717 34645 8751 34679
rect 8785 34645 8819 34679
rect 8853 34645 8887 34679
rect 8921 34645 8955 34679
rect 8989 34645 9023 34679
rect 9057 34645 9091 34679
rect 9125 34645 9159 34679
rect 9193 34645 9227 34679
rect 9261 34645 9295 34679
rect 9329 34645 9363 34679
rect 9397 34645 9431 34679
rect 9465 34645 9499 34679
rect 9533 34645 9567 34679
rect 9601 34645 9635 34679
rect 9669 34645 9703 34679
rect 9737 34645 9771 34679
rect 9805 34645 9839 34679
rect 9873 34645 9907 34679
rect 9941 34645 9975 34679
rect 10009 34645 10043 34679
rect 10077 34645 10111 34679
rect 10145 34645 10179 34679
rect 10213 34645 10247 34679
rect 10281 34645 10315 34679
rect 10349 34645 10383 34679
rect 10417 34645 10451 34679
rect 10485 34645 10519 34679
rect 10553 34645 10587 34679
rect 10621 34645 10655 34679
rect 10689 34645 10723 34679
rect 10757 34645 10791 34679
rect 10825 34645 10859 34679
rect 10893 34645 10927 34679
rect 10961 34645 10995 34679
rect 11029 34645 11063 34679
rect 11097 34645 11131 34679
rect 11165 34645 11199 34679
rect 11233 34645 11267 34679
rect 11301 34645 11335 34679
rect 11369 34645 11403 34679
rect 11437 34645 11471 34679
rect 11505 34645 11539 34679
rect 11573 34645 11607 34679
rect 11641 34645 11675 34679
rect 11709 34645 11743 34679
rect 11777 34645 11811 34679
rect 11845 34645 11879 34679
rect 11913 34645 11947 34679
rect 11981 34645 12015 34679
rect 12049 34645 12083 34679
rect 12117 34645 12151 34679
rect 12185 34645 12219 34679
rect 12253 34645 12287 34679
rect 12321 34645 12355 34679
rect 12389 34645 12423 34679
rect 12457 34645 12491 34679
rect 12525 34645 12559 34679
rect 12593 34645 12627 34679
rect 12661 34645 12695 34679
rect 12729 34645 12763 34679
rect 12797 34645 12831 34679
rect 12865 34645 12899 34679
rect 12933 34645 12967 34679
rect 13001 34645 13035 34679
rect 13069 34645 13103 34679
rect 13137 34645 13171 34679
rect 13205 34645 13239 34679
rect 13273 34645 13307 34679
rect 13341 34645 13375 34679
rect 13409 34645 13443 34679
rect 13477 34645 13511 34679
rect 13545 34645 13579 34679
rect 13613 34645 13647 34679
rect 13681 34645 13715 34679
rect 1161 34428 1195 34462
rect 1161 34360 1195 34394
rect 1161 34292 1195 34326
rect 1161 34224 1195 34258
rect 1161 34156 1195 34190
rect 1161 34088 1195 34122
rect 1161 34020 1195 34054
rect 1161 33952 1195 33986
rect 1161 33884 1195 33918
rect 1161 33816 1195 33850
rect 1161 33748 1195 33782
rect 1161 33680 1195 33714
rect 1161 33612 1195 33646
rect 1161 33544 1195 33578
rect 1161 33476 1195 33510
rect 1161 33408 1195 33442
rect 1161 33340 1195 33374
rect 1161 33272 1195 33306
rect 1161 33204 1195 33238
rect 1161 33136 1195 33170
rect 1161 33068 1195 33102
rect 1161 33000 1195 33034
rect 1161 32932 1195 32966
rect 1161 32864 1195 32898
rect 1161 32796 1195 32830
rect 1161 32728 1195 32762
rect 1161 32660 1195 32694
rect 1161 32592 1195 32626
rect 1161 32524 1195 32558
rect 1161 32456 1195 32490
rect 1161 32388 1195 32422
rect 1161 32320 1195 32354
rect 1161 32252 1195 32286
rect 1161 32184 1195 32218
rect 1161 32116 1195 32150
rect 1161 32048 1195 32082
rect 1161 31980 1195 32014
rect 1161 31912 1195 31946
rect 1161 31844 1195 31878
rect 1161 31776 1195 31810
rect 1161 31708 1195 31742
rect 1161 31640 1195 31674
rect 1161 31572 1195 31606
rect 1161 31504 1195 31538
rect 1161 31436 1195 31470
rect 1161 31368 1195 31402
rect 1161 31300 1195 31334
rect 1161 31232 1195 31266
rect 1161 31164 1195 31198
rect 1161 31096 1195 31130
rect 1161 31028 1195 31062
rect 1161 30960 1195 30994
rect 1161 30892 1195 30926
rect 1161 30824 1195 30858
rect 1161 30756 1195 30790
rect 1161 30688 1195 30722
rect 1161 30620 1195 30654
rect 1161 30552 1195 30586
rect 1161 30484 1195 30518
rect 1161 30416 1195 30450
rect 1161 30348 1195 30382
rect 1161 30280 1195 30314
rect 1161 30212 1195 30246
rect 1161 30144 1195 30178
rect 1161 30076 1195 30110
rect 1161 30008 1195 30042
rect 1161 29940 1195 29974
rect 1161 29872 1195 29906
rect 1161 29804 1195 29838
rect 1161 29736 1195 29770
rect 1161 29668 1195 29702
rect 1161 29600 1195 29634
rect 1161 29532 1195 29566
rect 1161 29464 1195 29498
rect 1161 29396 1195 29430
rect 1161 29328 1195 29362
rect 1161 29260 1195 29294
rect 1161 29192 1195 29226
rect 1161 29124 1195 29158
rect 1161 29056 1195 29090
rect 1161 28988 1195 29022
rect 1161 28920 1195 28954
rect 13809 34423 13843 34457
rect 13809 34355 13843 34389
rect 13809 34287 13843 34321
rect 13809 34219 13843 34253
rect 13809 34151 13843 34185
rect 13809 34083 13843 34117
rect 13809 34015 13843 34049
rect 13809 33947 13843 33981
rect 13809 33879 13843 33913
rect 13809 33811 13843 33845
rect 13809 33743 13843 33777
rect 13809 33675 13843 33709
rect 13809 33607 13843 33641
rect 13809 33539 13843 33573
rect 13809 33471 13843 33505
rect 13809 33403 13843 33437
rect 13809 33335 13843 33369
rect 13809 33267 13843 33301
rect 13809 33199 13843 33233
rect 13809 33131 13843 33165
rect 13809 33063 13843 33097
rect 13809 32995 13843 33029
rect 13809 32927 13843 32961
rect 13809 32859 13843 32893
rect 13809 32791 13843 32825
rect 13809 32723 13843 32757
rect 13809 32655 13843 32689
rect 13809 32587 13843 32621
rect 13809 32519 13843 32553
rect 13809 32451 13843 32485
rect 13809 32383 13843 32417
rect 13809 32315 13843 32349
rect 13809 32247 13843 32281
rect 13809 32179 13843 32213
rect 13809 32111 13843 32145
rect 13809 32043 13843 32077
rect 13809 31975 13843 32009
rect 13809 31907 13843 31941
rect 13809 31839 13843 31873
rect 13809 31771 13843 31805
rect 13809 31703 13843 31737
rect 13809 31635 13843 31669
rect 13809 31567 13843 31601
rect 13809 31499 13843 31533
rect 13809 31431 13843 31465
rect 13809 31363 13843 31397
rect 13809 31295 13843 31329
rect 13809 31227 13843 31261
rect 13809 31159 13843 31193
rect 13809 31091 13843 31125
rect 13809 31023 13843 31057
rect 13809 30955 13843 30989
rect 13809 30887 13843 30921
rect 13809 30819 13843 30853
rect 13809 30751 13843 30785
rect 13809 30683 13843 30717
rect 13809 30615 13843 30649
rect 13809 30547 13843 30581
rect 13809 30479 13843 30513
rect 13809 30411 13843 30445
rect 13809 30343 13843 30377
rect 13809 30275 13843 30309
rect 13809 30207 13843 30241
rect 13809 30139 13843 30173
rect 13809 30071 13843 30105
rect 13809 30003 13843 30037
rect 13809 29935 13843 29969
rect 13809 29867 13843 29901
rect 13809 29799 13843 29833
rect 13809 29731 13843 29765
rect 13809 29663 13843 29697
rect 13809 29595 13843 29629
rect 13809 29527 13843 29561
rect 13809 29459 13843 29493
rect 13809 29391 13843 29425
rect 13809 29323 13843 29357
rect 13809 29255 13843 29289
rect 13809 29187 13843 29221
rect 13809 29119 13843 29153
rect 13809 29051 13843 29085
rect 13809 28983 13843 29017
rect 13809 28915 13843 28949
rect 1161 28852 1195 28886
rect 1161 28784 1195 28818
rect 1161 28716 1195 28750
rect 1161 28648 1195 28682
rect 1161 28580 1195 28614
rect 1161 28512 1195 28546
rect 1161 28444 1195 28478
rect 1161 28376 1195 28410
rect 1161 28308 1195 28342
rect 1161 28240 1195 28274
rect 1161 28172 1195 28206
rect 1161 28104 1195 28138
rect 1161 28036 1195 28070
rect 1161 27968 1195 28002
rect 1161 27900 1195 27934
rect 1161 27832 1195 27866
rect 1161 27764 1195 27798
rect 1161 27696 1195 27730
rect 1161 27628 1195 27662
rect 1161 27560 1195 27594
rect 1161 27492 1195 27526
rect 1161 27424 1195 27458
rect 1161 27356 1195 27390
rect 1161 27288 1195 27322
rect 1161 27220 1195 27254
rect 1161 27152 1195 27186
rect 1161 27084 1195 27118
rect 1161 27016 1195 27050
rect 13809 28847 13843 28881
rect 13809 28779 13843 28813
rect 13809 28711 13843 28745
rect 13809 28643 13843 28677
rect 13809 28575 13843 28609
rect 13809 28507 13843 28541
rect 13809 28439 13843 28473
rect 13809 28371 13843 28405
rect 13809 28303 13843 28337
rect 13809 28235 13843 28269
rect 13809 28167 13843 28201
rect 13809 28099 13843 28133
rect 13809 28031 13843 28065
rect 13809 27963 13843 27997
rect 13809 27895 13843 27929
rect 13809 27827 13843 27861
rect 13809 27759 13843 27793
rect 13809 27691 13843 27725
rect 13809 27623 13843 27657
rect 13809 27555 13843 27589
rect 13809 27487 13843 27521
rect 13809 27419 13843 27453
rect 13809 27351 13843 27385
rect 13809 27283 13843 27317
rect 13809 27215 13843 27249
rect 13809 27147 13843 27181
rect 13809 27079 13843 27113
rect 1161 26948 1195 26982
rect 1161 26880 1195 26914
rect 1161 26812 1195 26846
rect 1161 26744 1195 26778
rect 1161 26676 1195 26710
rect 1161 26608 1195 26642
rect 1161 26540 1195 26574
rect 1161 26472 1195 26506
rect 1161 26404 1195 26438
rect 1161 26336 1195 26370
rect 1161 26268 1195 26302
rect 1161 26200 1195 26234
rect 1161 26132 1195 26166
rect 1161 26064 1195 26098
rect 1161 25996 1195 26030
rect 1161 25928 1195 25962
rect 1161 25860 1195 25894
rect 1161 25792 1195 25826
rect 1161 25724 1195 25758
rect 1161 25656 1195 25690
rect 1161 25588 1195 25622
rect 1161 25520 1195 25554
rect 1161 25452 1195 25486
rect 1161 25384 1195 25418
rect 1161 25316 1195 25350
rect 1161 25248 1195 25282
rect 1161 25180 1195 25214
rect 1161 25112 1195 25146
rect 1161 25044 1195 25078
rect 1161 24976 1195 25010
rect 1161 24908 1195 24942
rect 1161 24840 1195 24874
rect 1161 24772 1195 24806
rect 1161 24704 1195 24738
rect 1161 24636 1195 24670
rect 1161 24568 1195 24602
rect 1161 24500 1195 24534
rect 1161 24432 1195 24466
rect 1161 24364 1195 24398
rect 1161 24296 1195 24330
rect 1161 24228 1195 24262
rect 1161 24160 1195 24194
rect 1161 24092 1195 24126
rect 1161 24024 1195 24058
rect 1161 23956 1195 23990
rect 1161 23888 1195 23922
rect 1161 23820 1195 23854
rect 1161 23752 1195 23786
rect 1161 23684 1195 23718
rect 1161 23616 1195 23650
rect 1161 23548 1195 23582
rect 1161 23480 1195 23514
rect 1161 23412 1195 23446
rect 1161 23344 1195 23378
rect 1161 23276 1195 23310
rect 1161 23208 1195 23242
rect 1161 23140 1195 23174
rect 1161 23072 1195 23106
rect 1161 23004 1195 23038
rect 1161 22936 1195 22970
rect 1161 22868 1195 22902
rect 1161 22800 1195 22834
rect 1161 22732 1195 22766
rect 1161 22664 1195 22698
rect 1161 22596 1195 22630
rect 1161 22528 1195 22562
rect 1161 22460 1195 22494
rect 1161 22392 1195 22426
rect 1161 22324 1195 22358
rect 1161 22256 1195 22290
rect 1161 22188 1195 22222
rect 1161 22120 1195 22154
rect 1161 22052 1195 22086
rect 1161 21984 1195 22018
rect 1161 21916 1195 21950
rect 1161 21848 1195 21882
rect 1161 21780 1195 21814
rect 1161 21712 1195 21746
rect 1161 21644 1195 21678
rect 1161 21576 1195 21610
rect 1161 21508 1195 21542
rect 1161 21440 1195 21474
rect 1161 21372 1195 21406
rect 1161 21304 1195 21338
rect 1161 21236 1195 21270
rect 1161 21168 1195 21202
rect 1161 21100 1195 21134
rect 1161 21032 1195 21066
rect 1161 20964 1195 20998
rect 1161 20896 1195 20930
rect 1161 20828 1195 20862
rect 1161 20760 1195 20794
rect 1161 20692 1195 20726
rect 1161 20624 1195 20658
rect 1161 20556 1195 20590
rect 1161 20488 1195 20522
rect 1161 20420 1195 20454
rect 1161 20352 1195 20386
rect 1161 20284 1195 20318
rect 1161 20216 1195 20250
rect 1161 20148 1195 20182
rect 1161 20080 1195 20114
rect 1161 20012 1195 20046
rect 1161 19944 1195 19978
rect 1161 19876 1195 19910
rect 1161 19808 1195 19842
rect 1161 19740 1195 19774
rect 1161 19672 1195 19706
rect 1161 19604 1195 19638
rect 1161 19536 1195 19570
rect 1161 19468 1195 19502
rect 1161 19400 1195 19434
rect 1161 19332 1195 19366
rect 1161 19264 1195 19298
rect 1161 19196 1195 19230
rect 1161 19128 1195 19162
rect 1161 19060 1195 19094
rect 1161 18992 1195 19026
rect 1161 18924 1195 18958
rect 1161 18856 1195 18890
rect 1161 18788 1195 18822
rect 1161 18720 1195 18754
rect 1161 18652 1195 18686
rect 1161 18584 1195 18618
rect 1161 18516 1195 18550
rect 1161 18448 1195 18482
rect 1161 18380 1195 18414
rect 1161 18312 1195 18346
rect 1161 18244 1195 18278
rect 1161 18176 1195 18210
rect 1161 18108 1195 18142
rect 1161 18040 1195 18074
rect 1161 17972 1195 18006
rect 1161 17904 1195 17938
rect 1161 17836 1195 17870
rect 1161 17768 1195 17802
rect 1161 17700 1195 17734
rect 1161 17632 1195 17666
rect 1161 17564 1195 17598
rect 1161 17496 1195 17530
rect 1161 17428 1195 17462
rect 1161 17360 1195 17394
rect 1161 17292 1195 17326
rect 1161 17224 1195 17258
rect 1161 17156 1195 17190
rect 1161 17088 1195 17122
rect 1161 17020 1195 17054
rect 1161 16952 1195 16986
rect 1161 16884 1195 16918
rect 1161 16816 1195 16850
rect 1161 16748 1195 16782
rect 1161 16680 1195 16714
rect 1161 16612 1195 16646
rect 1161 16544 1195 16578
rect 1161 16476 1195 16510
rect 1161 16408 1195 16442
rect 1161 16340 1195 16374
rect 1161 16272 1195 16306
rect 1161 16204 1195 16238
rect 1161 16136 1195 16170
rect 1161 16068 1195 16102
rect 1161 16000 1195 16034
rect 1161 15932 1195 15966
rect 1161 15864 1195 15898
rect 1161 15796 1195 15830
rect 1161 15728 1195 15762
rect 1161 15660 1195 15694
rect 1161 15592 1195 15626
rect 1161 15524 1195 15558
rect 1161 15456 1195 15490
rect 1161 15388 1195 15422
rect 13809 27011 13843 27045
rect 13809 26943 13843 26977
rect 13809 26875 13843 26909
rect 13809 26807 13843 26841
rect 13809 26739 13843 26773
rect 13809 26671 13843 26705
rect 13809 26603 13843 26637
rect 13809 26535 13843 26569
rect 13809 26467 13843 26501
rect 13809 26399 13843 26433
rect 13809 26331 13843 26365
rect 13809 26263 13843 26297
rect 13809 26195 13843 26229
rect 13809 26127 13843 26161
rect 13809 26059 13843 26093
rect 13809 25991 13843 26025
rect 13809 25923 13843 25957
rect 13809 25855 13843 25889
rect 13809 25787 13843 25821
rect 13809 25719 13843 25753
rect 13809 25651 13843 25685
rect 13809 25583 13843 25617
rect 13809 25515 13843 25549
rect 13809 25447 13843 25481
rect 13809 25379 13843 25413
rect 13809 25311 13843 25345
rect 13809 25243 13843 25277
rect 13809 25175 13843 25209
rect 13809 25107 13843 25141
rect 13809 25039 13843 25073
rect 13809 24971 13843 25005
rect 13809 24903 13843 24937
rect 13809 24835 13843 24869
rect 13809 24767 13843 24801
rect 13809 24699 13843 24733
rect 13809 24631 13843 24665
rect 13809 24563 13843 24597
rect 13809 24495 13843 24529
rect 13809 24427 13843 24461
rect 13809 24359 13843 24393
rect 13809 24291 13843 24325
rect 13809 24223 13843 24257
rect 13809 24155 13843 24189
rect 13809 24087 13843 24121
rect 13809 24019 13843 24053
rect 13809 23951 13843 23985
rect 13809 23883 13843 23917
rect 13809 23815 13843 23849
rect 13809 23747 13843 23781
rect 13809 23679 13843 23713
rect 13809 23611 13843 23645
rect 13809 23543 13843 23577
rect 13809 23475 13843 23509
rect 13809 23407 13843 23441
rect 13809 23339 13843 23373
rect 13809 23271 13843 23305
rect 13809 23203 13843 23237
rect 13809 23135 13843 23169
rect 13809 23067 13843 23101
rect 13809 22999 13843 23033
rect 13809 22931 13843 22965
rect 13809 22863 13843 22897
rect 13809 22795 13843 22829
rect 13809 22727 13843 22761
rect 13809 22659 13843 22693
rect 13809 22591 13843 22625
rect 13809 22523 13843 22557
rect 13809 22455 13843 22489
rect 13809 22387 13843 22421
rect 13809 22319 13843 22353
rect 13809 22251 13843 22285
rect 13809 22183 13843 22217
rect 13809 22115 13843 22149
rect 13809 22047 13843 22081
rect 13809 21979 13843 22013
rect 13809 21911 13843 21945
rect 13809 21843 13843 21877
rect 13809 21775 13843 21809
rect 13809 21707 13843 21741
rect 13809 21639 13843 21673
rect 13809 21571 13843 21605
rect 13809 21503 13843 21537
rect 13809 21435 13843 21469
rect 13809 21367 13843 21401
rect 13809 21299 13843 21333
rect 13809 21231 13843 21265
rect 13809 21163 13843 21197
rect 13809 21095 13843 21129
rect 13809 21027 13843 21061
rect 13809 20959 13843 20993
rect 13809 20891 13843 20925
rect 13809 20823 13843 20857
rect 13809 20755 13843 20789
rect 13809 20687 13843 20721
rect 13809 20619 13843 20653
rect 13809 20551 13843 20585
rect 13809 20483 13843 20517
rect 13809 20415 13843 20449
rect 13809 20347 13843 20381
rect 13809 20279 13843 20313
rect 13809 20211 13843 20245
rect 13809 20143 13843 20177
rect 13809 20075 13843 20109
rect 13809 20007 13843 20041
rect 13809 19939 13843 19973
rect 13809 19871 13843 19905
rect 13809 19803 13843 19837
rect 13809 19735 13843 19769
rect 13809 19667 13843 19701
rect 13809 19599 13843 19633
rect 13809 19531 13843 19565
rect 13809 19463 13843 19497
rect 13809 19395 13843 19429
rect 13809 19327 13843 19361
rect 13809 19259 13843 19293
rect 13809 19191 13843 19225
rect 13809 19123 13843 19157
rect 13809 19055 13843 19089
rect 13809 18987 13843 19021
rect 13809 18919 13843 18953
rect 13809 18851 13843 18885
rect 13809 18783 13843 18817
rect 13809 18715 13843 18749
rect 13809 18647 13843 18681
rect 13809 18579 13843 18613
rect 13809 18511 13843 18545
rect 13809 18443 13843 18477
rect 13809 18375 13843 18409
rect 13809 18307 13843 18341
rect 13809 18239 13843 18273
rect 13809 18171 13843 18205
rect 13809 18103 13843 18137
rect 13809 18035 13843 18069
rect 13809 17967 13843 18001
rect 13809 17899 13843 17933
rect 13809 17831 13843 17865
rect 13809 17763 13843 17797
rect 13809 17695 13843 17729
rect 13809 17627 13843 17661
rect 13809 17559 13843 17593
rect 13809 17491 13843 17525
rect 13809 17423 13843 17457
rect 13809 17355 13843 17389
rect 13809 17287 13843 17321
rect 13809 17219 13843 17253
rect 13809 17151 13843 17185
rect 13809 17083 13843 17117
rect 13809 17015 13843 17049
rect 13809 16947 13843 16981
rect 13809 16879 13843 16913
rect 13809 16811 13843 16845
rect 13809 16743 13843 16777
rect 13809 16675 13843 16709
rect 13809 16607 13843 16641
rect 13809 16539 13843 16573
rect 13809 16471 13843 16505
rect 13809 16403 13843 16437
rect 13809 16335 13843 16369
rect 13809 16267 13843 16301
rect 13809 16199 13843 16233
rect 13809 16131 13843 16165
rect 13809 16063 13843 16097
rect 13809 15995 13843 16029
rect 13809 15927 13843 15961
rect 13809 15859 13843 15893
rect 13809 15791 13843 15825
rect 13809 15723 13843 15757
rect 13809 15655 13843 15689
rect 13809 15587 13843 15621
rect 13809 15519 13843 15553
rect 13809 15451 13843 15485
rect 13809 15383 13843 15417
rect 1302 15244 1336 15278
rect 1370 15244 1404 15278
rect 1438 15244 1472 15278
rect 1506 15244 1540 15278
rect 1574 15244 1608 15278
rect 1642 15244 1676 15278
rect 1710 15244 1744 15278
rect 1778 15244 1812 15278
rect 1846 15244 1880 15278
rect 1914 15244 1948 15278
rect 1982 15244 2016 15278
rect 2050 15244 2084 15278
rect 2118 15244 2152 15278
rect 2186 15244 2220 15278
rect 2254 15244 2288 15278
rect 2322 15244 2356 15278
rect 2390 15244 2424 15278
rect 2458 15244 2492 15278
rect 2526 15244 2560 15278
rect 2594 15244 2628 15278
rect 2662 15244 2696 15278
rect 2730 15244 2764 15278
rect 2798 15244 2832 15278
rect 2866 15244 2900 15278
rect 2934 15244 2968 15278
rect 3002 15244 3036 15278
rect 3070 15244 3104 15278
rect 3138 15244 3172 15278
rect 3206 15244 3240 15278
rect 3274 15244 3308 15278
rect 3342 15244 3376 15278
rect 3410 15244 3444 15278
rect 3478 15244 3512 15278
rect 3546 15244 3580 15278
rect 3614 15244 3648 15278
rect 3682 15244 3716 15278
rect 3750 15244 3784 15278
rect 3818 15244 3852 15278
rect 3886 15244 3920 15278
rect 3954 15244 3988 15278
rect 4022 15244 4056 15278
rect 4090 15244 4124 15278
rect 4158 15244 4192 15278
rect 4226 15244 4260 15278
rect 4294 15244 4328 15278
rect 4362 15244 4396 15278
rect 4430 15244 4464 15278
rect 4498 15244 4532 15278
rect 4566 15244 4600 15278
rect 4634 15244 4668 15278
rect 4702 15244 4736 15278
rect 4770 15244 4804 15278
rect 4838 15244 4872 15278
rect 4906 15244 4940 15278
rect 4974 15244 5008 15278
rect 5042 15244 5076 15278
rect 5110 15244 5144 15278
rect 5178 15244 5212 15278
rect 5246 15244 5280 15278
rect 5314 15244 5348 15278
rect 5382 15244 5416 15278
rect 5450 15244 5484 15278
rect 5518 15244 5552 15278
rect 5586 15244 5620 15278
rect 5654 15244 5688 15278
rect 5722 15244 5756 15278
rect 5790 15244 5824 15278
rect 5858 15244 5892 15278
rect 5926 15244 5960 15278
rect 5994 15244 6028 15278
rect 6062 15244 6096 15278
rect 6130 15244 6164 15278
rect 6198 15244 6232 15278
rect 6266 15244 6300 15278
rect 6334 15244 6368 15278
rect 6402 15244 6436 15278
rect 6470 15244 6504 15278
rect 6538 15244 6572 15278
rect 6606 15244 6640 15278
rect 6674 15244 6708 15278
rect 6742 15244 6776 15278
rect 6810 15244 6844 15278
rect 6878 15244 6912 15278
rect 6946 15244 6980 15278
rect 7014 15244 7048 15278
rect 7082 15244 7116 15278
rect 7150 15244 7184 15278
rect 7218 15244 7252 15278
rect 7286 15244 7320 15278
rect 7354 15244 7388 15278
rect 7422 15244 7456 15278
rect 7490 15244 7524 15278
rect 7558 15244 7592 15278
rect 7626 15244 7660 15278
rect 7694 15244 7728 15278
rect 7762 15244 7796 15278
rect 7830 15244 7864 15278
rect 7898 15244 7932 15278
rect 7966 15244 8000 15278
rect 8034 15244 8068 15278
rect 8102 15244 8136 15278
rect 8170 15244 8204 15278
rect 8238 15244 8272 15278
rect 8306 15244 8340 15278
rect 8374 15244 8408 15278
rect 8442 15244 8476 15278
rect 8510 15244 8544 15278
rect 8578 15244 8612 15278
rect 8646 15244 8680 15278
rect 8714 15244 8748 15278
rect 8782 15244 8816 15278
rect 8850 15244 8884 15278
rect 8918 15244 8952 15278
rect 8986 15244 9020 15278
rect 9054 15244 9088 15278
rect 9122 15244 9156 15278
rect 9190 15244 9224 15278
rect 9258 15244 9292 15278
rect 9326 15244 9360 15278
rect 9394 15244 9428 15278
rect 9462 15244 9496 15278
rect 9530 15244 9564 15278
rect 9598 15244 9632 15278
rect 9666 15244 9700 15278
rect 9734 15244 9768 15278
rect 9802 15244 9836 15278
rect 9870 15244 9904 15278
rect 9938 15244 9972 15278
rect 10006 15244 10040 15278
rect 10074 15244 10108 15278
rect 10142 15244 10176 15278
rect 10210 15244 10244 15278
rect 10278 15244 10312 15278
rect 10346 15244 10380 15278
rect 10414 15244 10448 15278
rect 10482 15244 10516 15278
rect 10550 15244 10584 15278
rect 10618 15244 10652 15278
rect 10686 15244 10720 15278
rect 10754 15244 10788 15278
rect 10822 15244 10856 15278
rect 10890 15244 10924 15278
rect 10958 15244 10992 15278
rect 11026 15244 11060 15278
rect 11094 15244 11128 15278
rect 11162 15244 11196 15278
rect 11230 15244 11264 15278
rect 11298 15244 11332 15278
rect 11366 15244 11400 15278
rect 11434 15244 11468 15278
rect 11502 15244 11536 15278
rect 11570 15244 11604 15278
rect 11638 15244 11672 15278
rect 11706 15244 11740 15278
rect 11774 15244 11808 15278
rect 11842 15244 11876 15278
rect 11910 15244 11944 15278
rect 11978 15244 12012 15278
rect 12046 15244 12080 15278
rect 12114 15244 12148 15278
rect 12182 15244 12216 15278
rect 12250 15244 12284 15278
rect 12318 15244 12352 15278
rect 12386 15244 12420 15278
rect 12454 15244 12488 15278
rect 12522 15244 12556 15278
rect 12590 15244 12624 15278
rect 12658 15244 12692 15278
rect 12726 15244 12760 15278
rect 12794 15244 12828 15278
rect 12862 15244 12896 15278
rect 12930 15244 12964 15278
rect 12998 15244 13032 15278
rect 13066 15244 13100 15278
rect 13134 15244 13168 15278
rect 13202 15244 13236 15278
rect 13270 15244 13304 15278
rect 13338 15244 13372 15278
rect 13406 15244 13440 15278
rect 13474 15244 13508 15278
rect 13542 15244 13576 15278
rect 13610 15244 13644 15278
rect 13678 15244 13712 15278
rect 14607 36192 14641 36226
rect 14607 36124 14641 36158
rect 14607 36056 14641 36090
rect 14607 35988 14641 36022
rect 14607 35920 14641 35954
rect 14607 35852 14641 35886
rect 14607 35784 14641 35818
rect 14607 35716 14641 35750
rect 14607 35648 14641 35682
rect 14607 35580 14641 35614
rect 14607 35512 14641 35546
rect 14607 35444 14641 35478
rect 14607 35376 14641 35410
rect 14607 35308 14641 35342
rect 14607 35240 14641 35274
rect 14607 35172 14641 35206
rect 14607 35104 14641 35138
rect 14607 35036 14641 35070
rect 14607 34968 14641 35002
rect 14607 34900 14641 34934
rect 14607 34832 14641 34866
rect 14607 34764 14641 34798
rect 14607 34696 14641 34730
rect 14607 34628 14641 34662
rect 14607 34560 14641 34594
rect 14607 34492 14641 34526
rect 14607 34424 14641 34458
rect 14607 34356 14641 34390
rect 14607 34288 14641 34322
rect 14607 34220 14641 34254
rect 14607 34152 14641 34186
rect 14607 34084 14641 34118
rect 14607 34016 14641 34050
rect 14607 33948 14641 33982
rect 14607 33880 14641 33914
rect 14607 33812 14641 33846
rect 14607 33744 14641 33778
rect 14607 33676 14641 33710
rect 14607 33608 14641 33642
rect 14607 33540 14641 33574
rect 14607 33472 14641 33506
rect 14607 33404 14641 33438
rect 14607 33336 14641 33370
rect 14607 33268 14641 33302
rect 14607 33200 14641 33234
rect 14607 33132 14641 33166
rect 14607 33064 14641 33098
rect 14607 32996 14641 33030
rect 14607 32928 14641 32962
rect 14607 32860 14641 32894
rect 14607 32792 14641 32826
rect 14607 32724 14641 32758
rect 14607 32656 14641 32690
rect 14607 32588 14641 32622
rect 14607 32520 14641 32554
rect 14607 32452 14641 32486
rect 14607 32384 14641 32418
rect 14607 32316 14641 32350
rect 14607 32248 14641 32282
rect 14607 32180 14641 32214
rect 14607 32112 14641 32146
rect 14607 32044 14641 32078
rect 14607 31976 14641 32010
rect 14607 31908 14641 31942
rect 14607 31840 14641 31874
rect 14607 31772 14641 31806
rect 14607 31704 14641 31738
rect 14607 31636 14641 31670
rect 14607 31568 14641 31602
rect 14607 31500 14641 31534
rect 14607 31432 14641 31466
rect 14607 31364 14641 31398
rect 14607 31296 14641 31330
rect 14607 31228 14641 31262
rect 14607 31160 14641 31194
rect 14607 31092 14641 31126
rect 14607 31024 14641 31058
rect 14607 30956 14641 30990
rect 14607 30888 14641 30922
rect 14607 30820 14641 30854
rect 14607 30752 14641 30786
rect 14607 30684 14641 30718
rect 14607 30616 14641 30650
rect 14607 30548 14641 30582
rect 14607 30480 14641 30514
rect 14607 30412 14641 30446
rect 14607 30344 14641 30378
rect 14607 30276 14641 30310
rect 14607 30208 14641 30242
rect 14607 30140 14641 30174
rect 14607 30072 14641 30106
rect 14607 30004 14641 30038
rect 14607 29936 14641 29970
rect 14607 29868 14641 29902
rect 14607 29800 14641 29834
rect 14607 29732 14641 29766
rect 14607 29664 14641 29698
rect 14607 29596 14641 29630
rect 14607 29528 14641 29562
rect 14607 29460 14641 29494
rect 14607 29392 14641 29426
rect 14607 29324 14641 29358
rect 14607 29256 14641 29290
rect 14607 29188 14641 29222
rect 14607 29120 14641 29154
rect 14607 29052 14641 29086
rect 14607 28984 14641 29018
rect 14607 28916 14641 28950
rect 14607 28848 14641 28882
rect 14607 28780 14641 28814
rect 14607 28712 14641 28746
rect 14607 28644 14641 28678
rect 14607 28576 14641 28610
rect 14607 28508 14641 28542
rect 14607 28440 14641 28474
rect 14607 28372 14641 28406
rect 14607 28304 14641 28338
rect 14607 28236 14641 28270
rect 14607 28168 14641 28202
rect 14607 28100 14641 28134
rect 14607 28032 14641 28066
rect 14607 27964 14641 27998
rect 14607 27896 14641 27930
rect 14607 27828 14641 27862
rect 14607 27760 14641 27794
rect 14607 27692 14641 27726
rect 14607 27624 14641 27658
rect 14607 27556 14641 27590
rect 14607 27488 14641 27522
rect 14607 27420 14641 27454
rect 14607 27352 14641 27386
rect 14607 27284 14641 27318
rect 14607 27216 14641 27250
rect 14607 27148 14641 27182
rect 14607 27080 14641 27114
rect 14607 27012 14641 27046
rect 14607 26944 14641 26978
rect 14607 26876 14641 26910
rect 14607 26808 14641 26842
rect 14607 26740 14641 26774
rect 14607 26672 14641 26706
rect 14607 26604 14641 26638
rect 14607 26536 14641 26570
rect 14607 26468 14641 26502
rect 14607 26400 14641 26434
rect 14607 26332 14641 26366
rect 14607 26264 14641 26298
rect 14607 26196 14641 26230
rect 14607 26128 14641 26162
rect 14607 26060 14641 26094
rect 14607 25992 14641 26026
rect 14607 25924 14641 25958
rect 14607 25856 14641 25890
rect 14607 25788 14641 25822
rect 14607 25720 14641 25754
rect 14607 25652 14641 25686
rect 14607 25584 14641 25618
rect 14607 25516 14641 25550
rect 14607 25448 14641 25482
rect 14607 25380 14641 25414
rect 14607 25312 14641 25346
rect 14607 25244 14641 25278
rect 14607 25176 14641 25210
rect 14607 25108 14641 25142
rect 14607 25040 14641 25074
rect 14607 24972 14641 25006
rect 14607 24904 14641 24938
rect 14607 24836 14641 24870
rect 14607 24768 14641 24802
rect 14607 24700 14641 24734
rect 14607 24632 14641 24666
rect 14607 24564 14641 24598
rect 14607 24496 14641 24530
rect 14607 24428 14641 24462
rect 14607 24360 14641 24394
rect 14607 24292 14641 24326
rect 14607 24224 14641 24258
rect 14607 24156 14641 24190
rect 14607 24088 14641 24122
rect 14607 24020 14641 24054
rect 14607 23952 14641 23986
rect 14607 23884 14641 23918
rect 14607 23816 14641 23850
rect 14607 23748 14641 23782
rect 14607 23680 14641 23714
rect 14607 23612 14641 23646
rect 14607 23544 14641 23578
rect 14607 23476 14641 23510
rect 14607 23408 14641 23442
rect 14607 23340 14641 23374
rect 14607 23272 14641 23306
rect 14607 23204 14641 23238
rect 14607 23136 14641 23170
rect 14607 23068 14641 23102
rect 14607 23000 14641 23034
rect 14607 22932 14641 22966
rect 14607 22864 14641 22898
rect 14607 22796 14641 22830
rect 14607 22728 14641 22762
rect 14607 22660 14641 22694
rect 14607 22592 14641 22626
rect 14607 22524 14641 22558
rect 14607 22456 14641 22490
rect 14607 22388 14641 22422
rect 14607 22320 14641 22354
rect 14607 22252 14641 22286
rect 14607 22184 14641 22218
rect 14607 22116 14641 22150
rect 14607 22048 14641 22082
rect 14607 21980 14641 22014
rect 14607 21912 14641 21946
rect 14607 21844 14641 21878
rect 14607 21776 14641 21810
rect 14607 21708 14641 21742
rect 14607 21640 14641 21674
rect 14607 21572 14641 21606
rect 14607 21504 14641 21538
rect 14607 21436 14641 21470
rect 14607 21368 14641 21402
rect 14607 21300 14641 21334
rect 14607 21232 14641 21266
rect 14607 21164 14641 21198
rect 14607 21096 14641 21130
rect 14607 21028 14641 21062
rect 14607 20960 14641 20994
rect 14607 20892 14641 20926
rect 14607 20824 14641 20858
rect 14607 20756 14641 20790
rect 14607 20688 14641 20722
rect 14607 20620 14641 20654
rect 14607 20552 14641 20586
rect 14607 20484 14641 20518
rect 14607 20416 14641 20450
rect 14607 20348 14641 20382
rect 14607 20280 14641 20314
rect 14607 20212 14641 20246
rect 14607 20144 14641 20178
rect 14607 20076 14641 20110
rect 14607 20008 14641 20042
rect 14607 19940 14641 19974
rect 14607 19872 14641 19906
rect 14607 19804 14641 19838
rect 14607 19736 14641 19770
rect 14607 19668 14641 19702
rect 14607 19600 14641 19634
rect 14607 19532 14641 19566
rect 14607 19464 14641 19498
rect 14607 19396 14641 19430
rect 14607 19328 14641 19362
rect 14607 19260 14641 19294
rect 14607 19192 14641 19226
rect 14607 19124 14641 19158
rect 14607 19056 14641 19090
rect 14607 18988 14641 19022
rect 14607 18920 14641 18954
rect 14607 18852 14641 18886
rect 14607 18784 14641 18818
rect 14607 18716 14641 18750
rect 14607 18648 14641 18682
rect 14607 18580 14641 18614
rect 14607 18512 14641 18546
rect 14607 18444 14641 18478
rect 14607 18376 14641 18410
rect 14607 18308 14641 18342
rect 14607 18240 14641 18274
rect 14607 18172 14641 18206
rect 14607 18104 14641 18138
rect 14607 18036 14641 18070
rect 14607 17968 14641 18002
rect 14607 17900 14641 17934
rect 14607 17832 14641 17866
rect 14607 17764 14641 17798
rect 14607 17696 14641 17730
rect 14607 17628 14641 17662
rect 14607 17560 14641 17594
rect 14607 17492 14641 17526
rect 14607 17424 14641 17458
rect 14607 17356 14641 17390
rect 14607 17288 14641 17322
rect 14607 17220 14641 17254
rect 14607 17152 14641 17186
rect 14607 17084 14641 17118
rect 14607 17016 14641 17050
rect 14607 16948 14641 16982
rect 14607 16880 14641 16914
rect 14607 16812 14641 16846
rect 14607 16744 14641 16778
rect 14607 16676 14641 16710
rect 14607 16608 14641 16642
rect 14607 16540 14641 16574
rect 14607 16472 14641 16506
rect 14607 16404 14641 16438
rect 14607 16336 14641 16370
rect 14607 16268 14641 16302
rect 14607 16200 14641 16234
rect 14607 16132 14641 16166
rect 14607 16064 14641 16098
rect 14607 15996 14641 16030
rect 14607 15928 14641 15962
rect 14607 15860 14641 15894
rect 14607 15792 14641 15826
rect 14607 15724 14641 15758
rect 14607 15656 14641 15690
rect 14607 15588 14641 15622
rect 14607 15520 14641 15554
rect 14607 15452 14641 15486
rect 14607 15384 14641 15418
rect 14607 15316 14641 15350
rect 14607 15248 14641 15282
rect 14607 15180 14641 15214
rect 14607 15112 14641 15146
rect 14607 15044 14641 15078
rect 14607 14976 14641 15010
rect 14607 14908 14641 14942
rect 14607 14840 14641 14874
rect 14607 14772 14641 14806
rect 14607 14704 14641 14738
rect 312 14630 346 14664
rect 312 14562 346 14596
rect 14607 14636 14641 14670
rect 14607 14568 14641 14602
rect 476 14417 510 14451
rect 544 14417 578 14451
rect 612 14417 646 14451
rect 680 14417 714 14451
rect 748 14417 782 14451
rect 816 14417 850 14451
rect 884 14417 918 14451
rect 952 14417 986 14451
rect 1020 14417 1054 14451
rect 1088 14417 1122 14451
rect 1156 14417 1190 14451
rect 1224 14417 1258 14451
rect 1292 14417 1326 14451
rect 1360 14417 1394 14451
rect 1428 14417 1462 14451
rect 1496 14417 1530 14451
rect 1564 14417 1598 14451
rect 1632 14417 1666 14451
rect 1700 14417 1734 14451
rect 1768 14417 1802 14451
rect 1836 14417 1870 14451
rect 1904 14417 1938 14451
rect 1972 14417 2006 14451
rect 2040 14417 2074 14451
rect 2108 14417 2142 14451
rect 2176 14417 2210 14451
rect 2244 14417 2278 14451
rect 2312 14417 2346 14451
rect 2380 14417 2414 14451
rect 2448 14417 2482 14451
rect 2516 14417 2550 14451
rect 2584 14417 2618 14451
rect 2652 14417 2686 14451
rect 2720 14417 2754 14451
rect 2788 14417 2822 14451
rect 2856 14417 2890 14451
rect 2924 14417 2958 14451
rect 2992 14417 3026 14451
rect 3060 14417 3094 14451
rect 3128 14417 3162 14451
rect 3196 14417 3230 14451
rect 3264 14417 3298 14451
rect 3332 14417 3366 14451
rect 3400 14417 3434 14451
rect 3468 14417 3502 14451
rect 3536 14417 3570 14451
rect 3604 14417 3638 14451
rect 3672 14417 3706 14451
rect 3740 14417 3774 14451
rect 3808 14417 3842 14451
rect 3876 14417 3910 14451
rect 3944 14417 3978 14451
rect 4012 14417 4046 14451
rect 4080 14417 4114 14451
rect 4148 14417 4182 14451
rect 4216 14417 4250 14451
rect 4284 14417 4318 14451
rect 4352 14417 4386 14451
rect 4420 14417 4454 14451
rect 4488 14417 4522 14451
rect 4556 14417 4590 14451
rect 4624 14417 4658 14451
rect 4692 14417 4726 14451
rect 4760 14417 4794 14451
rect 4828 14417 4862 14451
rect 4896 14417 4930 14451
rect 4964 14417 4998 14451
rect 5032 14417 5066 14451
rect 5100 14417 5134 14451
rect 5168 14417 5202 14451
rect 5236 14417 5270 14451
rect 5304 14417 5338 14451
rect 5372 14417 5406 14451
rect 5440 14417 5474 14451
rect 5508 14417 5542 14451
rect 5576 14417 5610 14451
rect 5644 14417 5678 14451
rect 5712 14417 5746 14451
rect 5780 14417 5814 14451
rect 5848 14417 5882 14451
rect 5916 14417 5950 14451
rect 5984 14417 6018 14451
rect 6052 14417 6086 14451
rect 6120 14417 6154 14451
rect 6188 14417 6222 14451
rect 6256 14417 6290 14451
rect 6324 14417 6358 14451
rect 6392 14417 6426 14451
rect 6460 14417 6494 14451
rect 6528 14417 6562 14451
rect 6596 14417 6630 14451
rect 6664 14417 6698 14451
rect 6732 14417 6766 14451
rect 6800 14417 6834 14451
rect 6868 14417 6902 14451
rect 6936 14417 6970 14451
rect 7004 14417 7038 14451
rect 7072 14417 7106 14451
rect 7140 14417 7174 14451
rect 7208 14417 7242 14451
rect 7276 14417 7310 14451
rect 7344 14417 7378 14451
rect 7412 14417 7446 14451
rect 7480 14417 7514 14451
rect 7548 14417 7582 14451
rect 7616 14417 7650 14451
rect 7684 14417 7718 14451
rect 7752 14417 7786 14451
rect 7820 14417 7854 14451
rect 7888 14417 7922 14451
rect 7956 14417 7990 14451
rect 8024 14417 8058 14451
rect 8092 14417 8126 14451
rect 8160 14417 8194 14451
rect 8228 14417 8262 14451
rect 8296 14417 8330 14451
rect 8364 14417 8398 14451
rect 8432 14417 8466 14451
rect 8500 14417 8534 14451
rect 8568 14417 8602 14451
rect 8636 14417 8670 14451
rect 8704 14417 8738 14451
rect 8772 14417 8806 14451
rect 8840 14417 8874 14451
rect 8908 14417 8942 14451
rect 8976 14417 9010 14451
rect 9044 14417 9078 14451
rect 9112 14417 9146 14451
rect 9180 14417 9214 14451
rect 9248 14417 9282 14451
rect 9316 14417 9350 14451
rect 9384 14417 9418 14451
rect 9452 14417 9486 14451
rect 9520 14417 9554 14451
rect 9588 14417 9622 14451
rect 9656 14417 9690 14451
rect 9724 14417 9758 14451
rect 9792 14417 9826 14451
rect 9860 14417 9894 14451
rect 9928 14417 9962 14451
rect 9996 14417 10030 14451
rect 10064 14417 10098 14451
rect 10132 14417 10166 14451
rect 10200 14417 10234 14451
rect 10268 14417 10302 14451
rect 10336 14417 10370 14451
rect 10404 14417 10438 14451
rect 10472 14417 10506 14451
rect 10540 14417 10574 14451
rect 10608 14417 10642 14451
rect 10676 14417 10710 14451
rect 10744 14417 10778 14451
rect 10812 14417 10846 14451
rect 10880 14417 10914 14451
rect 10948 14417 10982 14451
rect 11016 14417 11050 14451
rect 11084 14417 11118 14451
rect 11152 14417 11186 14451
rect 11220 14417 11254 14451
rect 11288 14417 11322 14451
rect 11356 14417 11390 14451
rect 11424 14417 11458 14451
rect 11492 14417 11526 14451
rect 11560 14417 11594 14451
rect 11628 14417 11662 14451
rect 11696 14417 11730 14451
rect 11764 14417 11798 14451
rect 11832 14417 11866 14451
rect 11900 14417 11934 14451
rect 11968 14417 12002 14451
rect 12036 14417 12070 14451
rect 12104 14417 12138 14451
rect 12172 14417 12206 14451
rect 12240 14417 12274 14451
rect 12308 14417 12342 14451
rect 12376 14417 12410 14451
rect 12444 14417 12478 14451
rect 12512 14417 12546 14451
rect 12580 14417 12614 14451
rect 12648 14417 12682 14451
rect 12716 14417 12750 14451
rect 12784 14417 12818 14451
rect 12852 14417 12886 14451
rect 12920 14417 12954 14451
rect 12988 14417 13022 14451
rect 13056 14417 13090 14451
rect 13124 14417 13158 14451
rect 13192 14417 13226 14451
rect 13260 14417 13294 14451
rect 13328 14417 13362 14451
rect 13396 14417 13430 14451
rect 13464 14417 13498 14451
rect 13532 14417 13566 14451
rect 13600 14417 13634 14451
rect 13668 14417 13702 14451
rect 13736 14417 13770 14451
rect 13804 14417 13838 14451
rect 13872 14417 13906 14451
rect 13940 14417 13974 14451
rect 14008 14417 14042 14451
rect 14076 14417 14110 14451
rect 14144 14417 14178 14451
rect 14212 14417 14246 14451
rect 14280 14417 14314 14451
rect 14348 14417 14382 14451
rect 14416 14417 14450 14451
rect 14484 14417 14518 14451
<< mvnsubdiffcont >>
rect 766 36143 800 36177
rect 834 36143 868 36177
rect 902 36143 936 36177
rect 970 36143 1004 36177
rect 1038 36143 1072 36177
rect 1106 36143 1140 36177
rect 1174 36143 1208 36177
rect 1242 36143 1276 36177
rect 1310 36143 1344 36177
rect 1378 36143 1412 36177
rect 1446 36143 1480 36177
rect 1514 36143 1548 36177
rect 1582 36143 1616 36177
rect 1650 36143 1684 36177
rect 1718 36143 1752 36177
rect 1786 36143 1820 36177
rect 1854 36143 1888 36177
rect 1922 36143 1956 36177
rect 1990 36143 2024 36177
rect 2058 36143 2092 36177
rect 2126 36143 2160 36177
rect 2194 36143 2228 36177
rect 2262 36143 2296 36177
rect 2330 36143 2364 36177
rect 2398 36143 2432 36177
rect 2466 36143 2500 36177
rect 2534 36143 2568 36177
rect 2602 36143 2636 36177
rect 2670 36143 2704 36177
rect 2738 36143 2772 36177
rect 2806 36143 2840 36177
rect 2874 36143 2908 36177
rect 2942 36143 2976 36177
rect 3010 36143 3044 36177
rect 3078 36143 3112 36177
rect 3146 36143 3180 36177
rect 3214 36143 3248 36177
rect 3282 36143 3316 36177
rect 3350 36143 3384 36177
rect 3418 36143 3452 36177
rect 3486 36143 3520 36177
rect 3554 36143 3588 36177
rect 3622 36143 3656 36177
rect 3690 36143 3724 36177
rect 3758 36143 3792 36177
rect 3826 36143 3860 36177
rect 3894 36143 3928 36177
rect 3962 36143 3996 36177
rect 4030 36143 4064 36177
rect 4098 36143 4132 36177
rect 4166 36143 4200 36177
rect 4234 36143 4268 36177
rect 4302 36143 4336 36177
rect 4370 36143 4404 36177
rect 4438 36143 4472 36177
rect 4506 36143 4540 36177
rect 4574 36143 4608 36177
rect 4642 36143 4676 36177
rect 4710 36143 4744 36177
rect 4778 36143 4812 36177
rect 4846 36143 4880 36177
rect 4914 36143 4948 36177
rect 4982 36143 5016 36177
rect 5050 36143 5084 36177
rect 5118 36143 5152 36177
rect 5186 36143 5220 36177
rect 5254 36143 5288 36177
rect 5322 36143 5356 36177
rect 5390 36143 5424 36177
rect 5458 36143 5492 36177
rect 5526 36143 5560 36177
rect 5594 36143 5628 36177
rect 5662 36143 5696 36177
rect 5730 36143 5764 36177
rect 5798 36143 5832 36177
rect 5866 36143 5900 36177
rect 5934 36143 5968 36177
rect 6002 36143 6036 36177
rect 6070 36143 6104 36177
rect 6138 36143 6172 36177
rect 6206 36143 6240 36177
rect 6274 36143 6308 36177
rect 6342 36143 6376 36177
rect 6410 36143 6444 36177
rect 6478 36143 6512 36177
rect 6546 36143 6580 36177
rect 6614 36143 6648 36177
rect 6682 36143 6716 36177
rect 6750 36143 6784 36177
rect 6818 36143 6852 36177
rect 6886 36143 6920 36177
rect 6954 36143 6988 36177
rect 7022 36143 7056 36177
rect 7090 36143 7124 36177
rect 7158 36143 7192 36177
rect 7226 36143 7260 36177
rect 7294 36143 7328 36177
rect 7362 36143 7396 36177
rect 7430 36143 7464 36177
rect 7498 36143 7532 36177
rect 7566 36143 7600 36177
rect 7634 36143 7668 36177
rect 7702 36143 7736 36177
rect 7770 36143 7804 36177
rect 7838 36143 7872 36177
rect 7906 36143 7940 36177
rect 7974 36143 8008 36177
rect 8042 36143 8076 36177
rect 8110 36143 8144 36177
rect 8178 36143 8212 36177
rect 8246 36143 8280 36177
rect 8314 36143 8348 36177
rect 8382 36143 8416 36177
rect 8450 36143 8484 36177
rect 8518 36143 8552 36177
rect 8586 36143 8620 36177
rect 8654 36143 8688 36177
rect 8722 36143 8756 36177
rect 8790 36143 8824 36177
rect 8858 36143 8892 36177
rect 8926 36143 8960 36177
rect 8994 36143 9028 36177
rect 9062 36143 9096 36177
rect 9130 36143 9164 36177
rect 9198 36143 9232 36177
rect 9266 36143 9300 36177
rect 9334 36143 9368 36177
rect 9402 36143 9436 36177
rect 9470 36143 9504 36177
rect 9538 36143 9572 36177
rect 9606 36143 9640 36177
rect 9674 36143 9708 36177
rect 9742 36143 9776 36177
rect 9810 36143 9844 36177
rect 9878 36143 9912 36177
rect 9946 36143 9980 36177
rect 10014 36143 10048 36177
rect 10082 36143 10116 36177
rect 10150 36143 10184 36177
rect 10218 36143 10252 36177
rect 10286 36143 10320 36177
rect 10354 36143 10388 36177
rect 10422 36143 10456 36177
rect 10490 36143 10524 36177
rect 10558 36143 10592 36177
rect 10626 36143 10660 36177
rect 10694 36143 10728 36177
rect 10762 36143 10796 36177
rect 10830 36143 10864 36177
rect 10898 36143 10932 36177
rect 10966 36143 11000 36177
rect 11034 36143 11068 36177
rect 11102 36143 11136 36177
rect 11170 36143 11204 36177
rect 11238 36143 11272 36177
rect 11306 36143 11340 36177
rect 11374 36143 11408 36177
rect 11442 36143 11476 36177
rect 11510 36143 11544 36177
rect 11578 36143 11612 36177
rect 11646 36143 11680 36177
rect 11714 36143 11748 36177
rect 11782 36143 11816 36177
rect 11850 36143 11884 36177
rect 11918 36143 11952 36177
rect 11986 36143 12020 36177
rect 12054 36143 12088 36177
rect 12122 36143 12156 36177
rect 12190 36143 12224 36177
rect 12258 36143 12292 36177
rect 12326 36143 12360 36177
rect 12394 36143 12428 36177
rect 12462 36143 12496 36177
rect 12530 36143 12564 36177
rect 12598 36143 12632 36177
rect 12666 36143 12700 36177
rect 12734 36143 12768 36177
rect 12802 36143 12836 36177
rect 12870 36143 12904 36177
rect 12938 36143 12972 36177
rect 13006 36143 13040 36177
rect 13074 36143 13108 36177
rect 13142 36143 13176 36177
rect 13210 36143 13244 36177
rect 13278 36143 13312 36177
rect 13346 36143 13380 36177
rect 13414 36143 13448 36177
rect 13482 36143 13516 36177
rect 13550 36143 13584 36177
rect 13618 36143 13652 36177
rect 13686 36143 13720 36177
rect 13754 36143 13788 36177
rect 13822 36143 13856 36177
rect 13890 36143 13924 36177
rect 13958 36143 13992 36177
rect 14026 36143 14060 36177
rect 14094 36143 14128 36177
rect 14162 36143 14196 36177
rect 632 36016 666 36050
rect 632 35948 666 35982
rect 632 35880 666 35914
rect 632 35812 666 35846
rect 632 35744 666 35778
rect 632 35676 666 35710
rect 632 35608 666 35642
rect 632 35540 666 35574
rect 632 35472 666 35506
rect 632 35404 666 35438
rect 632 35336 666 35370
rect 632 35268 666 35302
rect 632 35200 666 35234
rect 632 35132 666 35166
rect 632 35064 666 35098
rect 632 34996 666 35030
rect 632 34928 666 34962
rect 632 34860 666 34894
rect 632 34792 666 34826
rect 632 34724 666 34758
rect 14297 36016 14331 36050
rect 14297 35948 14331 35982
rect 14297 35880 14331 35914
rect 14297 35812 14331 35846
rect 14297 35744 14331 35778
rect 14297 35676 14331 35710
rect 14297 35608 14331 35642
rect 14297 35540 14331 35574
rect 14297 35472 14331 35506
rect 14297 35404 14331 35438
rect 14297 35336 14331 35370
rect 14297 35268 14331 35302
rect 14297 35200 14331 35234
rect 14297 35132 14331 35166
rect 14297 35064 14331 35098
rect 14297 34996 14331 35030
rect 14297 34928 14331 34962
rect 14297 34860 14331 34894
rect 14297 34792 14331 34826
rect 14297 34724 14331 34758
rect 632 34656 666 34690
rect 632 34588 666 34622
rect 632 34520 666 34554
rect 632 34452 666 34486
rect 632 34384 666 34418
rect 632 34316 666 34350
rect 632 34248 666 34282
rect 632 34180 666 34214
rect 632 34112 666 34146
rect 632 34044 666 34078
rect 632 33976 666 34010
rect 632 33908 666 33942
rect 632 33840 666 33874
rect 632 33772 666 33806
rect 632 33704 666 33738
rect 632 33636 666 33670
rect 632 33568 666 33602
rect 632 33500 666 33534
rect 632 33432 666 33466
rect 632 33364 666 33398
rect 632 33296 666 33330
rect 632 33228 666 33262
rect 632 33160 666 33194
rect 632 33092 666 33126
rect 632 33024 666 33058
rect 632 32956 666 32990
rect 632 32888 666 32922
rect 632 32820 666 32854
rect 632 32752 666 32786
rect 632 32684 666 32718
rect 632 32616 666 32650
rect 632 32548 666 32582
rect 632 32480 666 32514
rect 632 32412 666 32446
rect 632 32344 666 32378
rect 632 32276 666 32310
rect 632 32208 666 32242
rect 632 32140 666 32174
rect 632 32072 666 32106
rect 632 32004 666 32038
rect 632 31936 666 31970
rect 632 31868 666 31902
rect 632 31800 666 31834
rect 632 31732 666 31766
rect 632 31664 666 31698
rect 632 31596 666 31630
rect 632 31528 666 31562
rect 632 31460 666 31494
rect 632 31392 666 31426
rect 632 31324 666 31358
rect 632 31256 666 31290
rect 632 31188 666 31222
rect 632 31120 666 31154
rect 632 31052 666 31086
rect 632 30984 666 31018
rect 632 30916 666 30950
rect 632 30848 666 30882
rect 632 30780 666 30814
rect 632 30712 666 30746
rect 632 30644 666 30678
rect 632 30576 666 30610
rect 632 30508 666 30542
rect 632 30440 666 30474
rect 632 30372 666 30406
rect 632 30304 666 30338
rect 632 30236 666 30270
rect 632 30168 666 30202
rect 632 30100 666 30134
rect 632 30032 666 30066
rect 632 29964 666 29998
rect 632 29896 666 29930
rect 632 29828 666 29862
rect 632 29760 666 29794
rect 632 29692 666 29726
rect 632 29624 666 29658
rect 632 29556 666 29590
rect 632 29488 666 29522
rect 632 29420 666 29454
rect 632 29352 666 29386
rect 632 29284 666 29318
rect 632 29216 666 29250
rect 632 29148 666 29182
rect 632 29080 666 29114
rect 632 29012 666 29046
rect 632 28944 666 28978
rect 632 28876 666 28910
rect 632 28808 666 28842
rect 632 28740 666 28774
rect 632 28672 666 28706
rect 632 28604 666 28638
rect 632 28536 666 28570
rect 632 28468 666 28502
rect 632 28400 666 28434
rect 632 28332 666 28366
rect 632 28264 666 28298
rect 632 28196 666 28230
rect 632 28128 666 28162
rect 632 28060 666 28094
rect 632 27992 666 28026
rect 632 27924 666 27958
rect 632 27856 666 27890
rect 632 27788 666 27822
rect 632 27720 666 27754
rect 632 27652 666 27686
rect 632 27584 666 27618
rect 632 27516 666 27550
rect 632 27448 666 27482
rect 632 27380 666 27414
rect 632 27312 666 27346
rect 632 27244 666 27278
rect 632 27176 666 27210
rect 632 27108 666 27142
rect 632 27040 666 27074
rect 632 26972 666 27006
rect 632 26904 666 26938
rect 632 26836 666 26870
rect 632 26768 666 26802
rect 632 26700 666 26734
rect 632 26632 666 26666
rect 632 26564 666 26598
rect 632 26496 666 26530
rect 632 26428 666 26462
rect 632 26360 666 26394
rect 632 26292 666 26326
rect 632 26224 666 26258
rect 632 26156 666 26190
rect 632 26088 666 26122
rect 632 26020 666 26054
rect 632 25952 666 25986
rect 632 25884 666 25918
rect 632 25816 666 25850
rect 632 25748 666 25782
rect 632 25680 666 25714
rect 632 25612 666 25646
rect 632 25544 666 25578
rect 632 25476 666 25510
rect 632 25408 666 25442
rect 632 25340 666 25374
rect 632 25272 666 25306
rect 632 25204 666 25238
rect 632 25136 666 25170
rect 632 25068 666 25102
rect 632 25000 666 25034
rect 632 24932 666 24966
rect 632 24864 666 24898
rect 632 24796 666 24830
rect 632 24728 666 24762
rect 632 24660 666 24694
rect 632 24592 666 24626
rect 632 24524 666 24558
rect 632 24456 666 24490
rect 632 24388 666 24422
rect 632 24320 666 24354
rect 632 24252 666 24286
rect 632 24184 666 24218
rect 632 24116 666 24150
rect 632 24048 666 24082
rect 632 23980 666 24014
rect 632 23912 666 23946
rect 632 23844 666 23878
rect 632 23776 666 23810
rect 632 23708 666 23742
rect 632 23640 666 23674
rect 632 23572 666 23606
rect 632 23504 666 23538
rect 632 23436 666 23470
rect 632 23368 666 23402
rect 632 23300 666 23334
rect 632 23232 666 23266
rect 632 23164 666 23198
rect 632 23096 666 23130
rect 632 23028 666 23062
rect 632 22960 666 22994
rect 632 22892 666 22926
rect 632 22824 666 22858
rect 632 22756 666 22790
rect 632 22688 666 22722
rect 632 22620 666 22654
rect 632 22552 666 22586
rect 632 22484 666 22518
rect 632 22416 666 22450
rect 632 22348 666 22382
rect 632 22280 666 22314
rect 632 22212 666 22246
rect 632 22144 666 22178
rect 632 22076 666 22110
rect 632 22008 666 22042
rect 632 21940 666 21974
rect 632 21872 666 21906
rect 632 21804 666 21838
rect 632 21736 666 21770
rect 632 21668 666 21702
rect 632 21600 666 21634
rect 632 21532 666 21566
rect 632 21464 666 21498
rect 632 21396 666 21430
rect 632 21328 666 21362
rect 632 21260 666 21294
rect 632 21192 666 21226
rect 632 21124 666 21158
rect 632 21056 666 21090
rect 632 20988 666 21022
rect 632 20920 666 20954
rect 632 20852 666 20886
rect 632 20784 666 20818
rect 632 20716 666 20750
rect 632 20648 666 20682
rect 632 20580 666 20614
rect 632 20512 666 20546
rect 632 20444 666 20478
rect 632 20376 666 20410
rect 632 20308 666 20342
rect 632 20240 666 20274
rect 632 20172 666 20206
rect 632 20104 666 20138
rect 632 20036 666 20070
rect 632 19968 666 20002
rect 632 19900 666 19934
rect 632 19832 666 19866
rect 632 19764 666 19798
rect 632 19696 666 19730
rect 632 19628 666 19662
rect 632 19560 666 19594
rect 632 19492 666 19526
rect 632 19424 666 19458
rect 632 19356 666 19390
rect 632 19288 666 19322
rect 632 19220 666 19254
rect 632 19152 666 19186
rect 632 19084 666 19118
rect 632 19016 666 19050
rect 632 18948 666 18982
rect 632 18880 666 18914
rect 632 18812 666 18846
rect 632 18744 666 18778
rect 632 18676 666 18710
rect 632 18608 666 18642
rect 632 18540 666 18574
rect 632 18472 666 18506
rect 632 18404 666 18438
rect 632 18336 666 18370
rect 632 18268 666 18302
rect 632 18200 666 18234
rect 632 18132 666 18166
rect 632 18064 666 18098
rect 632 17996 666 18030
rect 632 17928 666 17962
rect 632 17860 666 17894
rect 632 17792 666 17826
rect 632 17724 666 17758
rect 632 17656 666 17690
rect 632 17588 666 17622
rect 632 17520 666 17554
rect 632 17452 666 17486
rect 632 17384 666 17418
rect 632 17316 666 17350
rect 632 17248 666 17282
rect 632 17180 666 17214
rect 632 17112 666 17146
rect 632 17044 666 17078
rect 632 16976 666 17010
rect 632 16908 666 16942
rect 632 16840 666 16874
rect 632 16772 666 16806
rect 632 16704 666 16738
rect 632 16636 666 16670
rect 632 16568 666 16602
rect 632 16500 666 16534
rect 632 16432 666 16466
rect 632 16364 666 16398
rect 632 16296 666 16330
rect 632 16228 666 16262
rect 632 16160 666 16194
rect 632 16092 666 16126
rect 632 16024 666 16058
rect 632 15956 666 15990
rect 632 15888 666 15922
rect 632 15820 666 15854
rect 632 15752 666 15786
rect 632 15684 666 15718
rect 632 15616 666 15650
rect 632 15548 666 15582
rect 632 15480 666 15514
rect 632 15412 666 15446
rect 632 15344 666 15378
rect 632 15276 666 15310
rect 632 15208 666 15242
rect 2119 28505 12897 28879
rect 1689 27504 2063 28422
rect 12953 27504 13327 28422
rect 2119 27047 12897 27421
rect 14297 34656 14331 34690
rect 14297 34588 14331 34622
rect 14297 34520 14331 34554
rect 14297 34452 14331 34486
rect 14297 34384 14331 34418
rect 14297 34316 14331 34350
rect 14297 34248 14331 34282
rect 14297 34180 14331 34214
rect 14297 34112 14331 34146
rect 14297 34044 14331 34078
rect 14297 33976 14331 34010
rect 14297 33908 14331 33942
rect 14297 33840 14331 33874
rect 14297 33772 14331 33806
rect 14297 33704 14331 33738
rect 14297 33636 14331 33670
rect 14297 33568 14331 33602
rect 14297 33500 14331 33534
rect 14297 33432 14331 33466
rect 14297 33364 14331 33398
rect 14297 33296 14331 33330
rect 14297 33228 14331 33262
rect 14297 33160 14331 33194
rect 14297 33092 14331 33126
rect 14297 33024 14331 33058
rect 14297 32956 14331 32990
rect 14297 32888 14331 32922
rect 14297 32820 14331 32854
rect 14297 32752 14331 32786
rect 14297 32684 14331 32718
rect 14297 32616 14331 32650
rect 14297 32548 14331 32582
rect 14297 32480 14331 32514
rect 14297 32412 14331 32446
rect 14297 32344 14331 32378
rect 14297 32276 14331 32310
rect 14297 32208 14331 32242
rect 14297 32140 14331 32174
rect 14297 32072 14331 32106
rect 14297 32004 14331 32038
rect 14297 31936 14331 31970
rect 14297 31868 14331 31902
rect 14297 31800 14331 31834
rect 14297 31732 14331 31766
rect 14297 31664 14331 31698
rect 14297 31596 14331 31630
rect 14297 31528 14331 31562
rect 14297 31460 14331 31494
rect 14297 31392 14331 31426
rect 14297 31324 14331 31358
rect 14297 31256 14331 31290
rect 14297 31188 14331 31222
rect 14297 31120 14331 31154
rect 14297 31052 14331 31086
rect 14297 30984 14331 31018
rect 14297 30916 14331 30950
rect 14297 30848 14331 30882
rect 14297 30780 14331 30814
rect 14297 30712 14331 30746
rect 14297 30644 14331 30678
rect 14297 30576 14331 30610
rect 14297 30508 14331 30542
rect 14297 30440 14331 30474
rect 14297 30372 14331 30406
rect 14297 30304 14331 30338
rect 14297 30236 14331 30270
rect 14297 30168 14331 30202
rect 14297 30100 14331 30134
rect 14297 30032 14331 30066
rect 14297 29964 14331 29998
rect 14297 29896 14331 29930
rect 14297 29828 14331 29862
rect 14297 29760 14331 29794
rect 14297 29692 14331 29726
rect 14297 29624 14331 29658
rect 14297 29556 14331 29590
rect 14297 29488 14331 29522
rect 14297 29420 14331 29454
rect 14297 29352 14331 29386
rect 14297 29284 14331 29318
rect 14297 29216 14331 29250
rect 14297 29148 14331 29182
rect 14297 29080 14331 29114
rect 14297 29012 14331 29046
rect 14297 28944 14331 28978
rect 14297 28876 14331 28910
rect 14297 28808 14331 28842
rect 14297 28740 14331 28774
rect 14297 28672 14331 28706
rect 14297 28604 14331 28638
rect 14297 28536 14331 28570
rect 14297 28468 14331 28502
rect 14297 28400 14331 28434
rect 14297 28332 14331 28366
rect 14297 28264 14331 28298
rect 14297 28196 14331 28230
rect 14297 28128 14331 28162
rect 14297 28060 14331 28094
rect 14297 27992 14331 28026
rect 14297 27924 14331 27958
rect 14297 27856 14331 27890
rect 14297 27788 14331 27822
rect 14297 27720 14331 27754
rect 14297 27652 14331 27686
rect 14297 27584 14331 27618
rect 14297 27516 14331 27550
rect 14297 27448 14331 27482
rect 14297 27380 14331 27414
rect 14297 27312 14331 27346
rect 14297 27244 14331 27278
rect 14297 27176 14331 27210
rect 14297 27108 14331 27142
rect 14297 27040 14331 27074
rect 14297 26972 14331 27006
rect 14297 26904 14331 26938
rect 14297 26836 14331 26870
rect 14297 26768 14331 26802
rect 14297 26700 14331 26734
rect 14297 26632 14331 26666
rect 14297 26564 14331 26598
rect 14297 26496 14331 26530
rect 14297 26428 14331 26462
rect 14297 26360 14331 26394
rect 14297 26292 14331 26326
rect 14297 26224 14331 26258
rect 14297 26156 14331 26190
rect 14297 26088 14331 26122
rect 14297 26020 14331 26054
rect 14297 25952 14331 25986
rect 14297 25884 14331 25918
rect 14297 25816 14331 25850
rect 14297 25748 14331 25782
rect 14297 25680 14331 25714
rect 14297 25612 14331 25646
rect 14297 25544 14331 25578
rect 14297 25476 14331 25510
rect 14297 25408 14331 25442
rect 14297 25340 14331 25374
rect 14297 25272 14331 25306
rect 14297 25204 14331 25238
rect 14297 25136 14331 25170
rect 14297 25068 14331 25102
rect 14297 25000 14331 25034
rect 14297 24932 14331 24966
rect 14297 24864 14331 24898
rect 14297 24796 14331 24830
rect 14297 24728 14331 24762
rect 14297 24660 14331 24694
rect 14297 24592 14331 24626
rect 14297 24524 14331 24558
rect 14297 24456 14331 24490
rect 14297 24388 14331 24422
rect 14297 24320 14331 24354
rect 14297 24252 14331 24286
rect 14297 24184 14331 24218
rect 14297 24116 14331 24150
rect 14297 24048 14331 24082
rect 14297 23980 14331 24014
rect 14297 23912 14331 23946
rect 14297 23844 14331 23878
rect 14297 23776 14331 23810
rect 14297 23708 14331 23742
rect 14297 23640 14331 23674
rect 14297 23572 14331 23606
rect 14297 23504 14331 23538
rect 14297 23436 14331 23470
rect 14297 23368 14331 23402
rect 14297 23300 14331 23334
rect 14297 23232 14331 23266
rect 14297 23164 14331 23198
rect 14297 23096 14331 23130
rect 14297 23028 14331 23062
rect 14297 22960 14331 22994
rect 14297 22892 14331 22926
rect 14297 22824 14331 22858
rect 14297 22756 14331 22790
rect 14297 22688 14331 22722
rect 14297 22620 14331 22654
rect 14297 22552 14331 22586
rect 14297 22484 14331 22518
rect 14297 22416 14331 22450
rect 14297 22348 14331 22382
rect 14297 22280 14331 22314
rect 14297 22212 14331 22246
rect 14297 22144 14331 22178
rect 14297 22076 14331 22110
rect 14297 22008 14331 22042
rect 14297 21940 14331 21974
rect 14297 21872 14331 21906
rect 14297 21804 14331 21838
rect 14297 21736 14331 21770
rect 14297 21668 14331 21702
rect 14297 21600 14331 21634
rect 14297 21532 14331 21566
rect 14297 21464 14331 21498
rect 14297 21396 14331 21430
rect 14297 21328 14331 21362
rect 14297 21260 14331 21294
rect 14297 21192 14331 21226
rect 14297 21124 14331 21158
rect 14297 21056 14331 21090
rect 14297 20988 14331 21022
rect 14297 20920 14331 20954
rect 14297 20852 14331 20886
rect 14297 20784 14331 20818
rect 14297 20716 14331 20750
rect 14297 20648 14331 20682
rect 14297 20580 14331 20614
rect 14297 20512 14331 20546
rect 14297 20444 14331 20478
rect 14297 20376 14331 20410
rect 14297 20308 14331 20342
rect 14297 20240 14331 20274
rect 14297 20172 14331 20206
rect 14297 20104 14331 20138
rect 14297 20036 14331 20070
rect 14297 19968 14331 20002
rect 14297 19900 14331 19934
rect 14297 19832 14331 19866
rect 14297 19764 14331 19798
rect 14297 19696 14331 19730
rect 14297 19628 14331 19662
rect 14297 19560 14331 19594
rect 14297 19492 14331 19526
rect 14297 19424 14331 19458
rect 14297 19356 14331 19390
rect 14297 19288 14331 19322
rect 14297 19220 14331 19254
rect 14297 19152 14331 19186
rect 14297 19084 14331 19118
rect 14297 19016 14331 19050
rect 14297 18948 14331 18982
rect 14297 18880 14331 18914
rect 14297 18812 14331 18846
rect 14297 18744 14331 18778
rect 14297 18676 14331 18710
rect 14297 18608 14331 18642
rect 14297 18540 14331 18574
rect 14297 18472 14331 18506
rect 14297 18404 14331 18438
rect 14297 18336 14331 18370
rect 14297 18268 14331 18302
rect 14297 18200 14331 18234
rect 14297 18132 14331 18166
rect 14297 18064 14331 18098
rect 14297 17996 14331 18030
rect 14297 17928 14331 17962
rect 14297 17860 14331 17894
rect 14297 17792 14331 17826
rect 14297 17724 14331 17758
rect 14297 17656 14331 17690
rect 14297 17588 14331 17622
rect 14297 17520 14331 17554
rect 14297 17452 14331 17486
rect 14297 17384 14331 17418
rect 14297 17316 14331 17350
rect 14297 17248 14331 17282
rect 14297 17180 14331 17214
rect 14297 17112 14331 17146
rect 14297 17044 14331 17078
rect 14297 16976 14331 17010
rect 14297 16908 14331 16942
rect 14297 16840 14331 16874
rect 14297 16772 14331 16806
rect 14297 16704 14331 16738
rect 14297 16636 14331 16670
rect 14297 16568 14331 16602
rect 14297 16500 14331 16534
rect 14297 16432 14331 16466
rect 14297 16364 14331 16398
rect 14297 16296 14331 16330
rect 14297 16228 14331 16262
rect 14297 16160 14331 16194
rect 14297 16092 14331 16126
rect 14297 16024 14331 16058
rect 14297 15956 14331 15990
rect 14297 15888 14331 15922
rect 14297 15820 14331 15854
rect 14297 15752 14331 15786
rect 14297 15684 14331 15718
rect 14297 15616 14331 15650
rect 14297 15548 14331 15582
rect 14297 15480 14331 15514
rect 14297 15412 14331 15446
rect 14297 15344 14331 15378
rect 14297 15276 14331 15310
rect 14297 15208 14331 15242
rect 632 15140 666 15174
rect 632 15072 666 15106
rect 632 15004 666 15038
rect 632 14936 666 14970
rect 632 14868 666 14902
rect 14297 15140 14331 15174
rect 14297 15072 14331 15106
rect 14297 15004 14331 15038
rect 14297 14936 14331 14970
rect 14297 14868 14331 14902
rect 766 14741 800 14775
rect 834 14741 868 14775
rect 902 14741 936 14775
rect 970 14741 1004 14775
rect 1038 14741 1072 14775
rect 1106 14741 1140 14775
rect 1174 14741 1208 14775
rect 1242 14741 1276 14775
rect 1310 14741 1344 14775
rect 1378 14741 1412 14775
rect 1446 14741 1480 14775
rect 1514 14741 1548 14775
rect 1582 14741 1616 14775
rect 1650 14741 1684 14775
rect 1718 14741 1752 14775
rect 1786 14741 1820 14775
rect 1854 14741 1888 14775
rect 1922 14741 1956 14775
rect 1990 14741 2024 14775
rect 2058 14741 2092 14775
rect 2126 14741 2160 14775
rect 2194 14741 2228 14775
rect 2262 14741 2296 14775
rect 2330 14741 2364 14775
rect 2398 14741 2432 14775
rect 2466 14741 2500 14775
rect 2534 14741 2568 14775
rect 2602 14741 2636 14775
rect 2670 14741 2704 14775
rect 2738 14741 2772 14775
rect 2806 14741 2840 14775
rect 2874 14741 2908 14775
rect 2942 14741 2976 14775
rect 3010 14741 3044 14775
rect 3078 14741 3112 14775
rect 3146 14741 3180 14775
rect 3214 14741 3248 14775
rect 3282 14741 3316 14775
rect 3350 14741 3384 14775
rect 3418 14741 3452 14775
rect 3486 14741 3520 14775
rect 3554 14741 3588 14775
rect 3622 14741 3656 14775
rect 3690 14741 3724 14775
rect 3758 14741 3792 14775
rect 3826 14741 3860 14775
rect 3894 14741 3928 14775
rect 3962 14741 3996 14775
rect 4030 14741 4064 14775
rect 4098 14741 4132 14775
rect 4166 14741 4200 14775
rect 4234 14741 4268 14775
rect 4302 14741 4336 14775
rect 4370 14741 4404 14775
rect 4438 14741 4472 14775
rect 4506 14741 4540 14775
rect 4574 14741 4608 14775
rect 4642 14741 4676 14775
rect 4710 14741 4744 14775
rect 4778 14741 4812 14775
rect 4846 14741 4880 14775
rect 4914 14741 4948 14775
rect 4982 14741 5016 14775
rect 5050 14741 5084 14775
rect 5118 14741 5152 14775
rect 5186 14741 5220 14775
rect 5254 14741 5288 14775
rect 5322 14741 5356 14775
rect 5390 14741 5424 14775
rect 5458 14741 5492 14775
rect 5526 14741 5560 14775
rect 5594 14741 5628 14775
rect 5662 14741 5696 14775
rect 5730 14741 5764 14775
rect 5798 14741 5832 14775
rect 5866 14741 5900 14775
rect 5934 14741 5968 14775
rect 6002 14741 6036 14775
rect 6070 14741 6104 14775
rect 6138 14741 6172 14775
rect 6206 14741 6240 14775
rect 6274 14741 6308 14775
rect 6342 14741 6376 14775
rect 6410 14741 6444 14775
rect 6478 14741 6512 14775
rect 6546 14741 6580 14775
rect 6614 14741 6648 14775
rect 6682 14741 6716 14775
rect 6750 14741 6784 14775
rect 6818 14741 6852 14775
rect 6886 14741 6920 14775
rect 6954 14741 6988 14775
rect 7022 14741 7056 14775
rect 7090 14741 7124 14775
rect 7158 14741 7192 14775
rect 7226 14741 7260 14775
rect 7294 14741 7328 14775
rect 7362 14741 7396 14775
rect 7430 14741 7464 14775
rect 7498 14741 7532 14775
rect 7566 14741 7600 14775
rect 7634 14741 7668 14775
rect 7702 14741 7736 14775
rect 7770 14741 7804 14775
rect 7838 14741 7872 14775
rect 7906 14741 7940 14775
rect 7974 14741 8008 14775
rect 8042 14741 8076 14775
rect 8110 14741 8144 14775
rect 8178 14741 8212 14775
rect 8246 14741 8280 14775
rect 8314 14741 8348 14775
rect 8382 14741 8416 14775
rect 8450 14741 8484 14775
rect 8518 14741 8552 14775
rect 8586 14741 8620 14775
rect 8654 14741 8688 14775
rect 8722 14741 8756 14775
rect 8790 14741 8824 14775
rect 8858 14741 8892 14775
rect 8926 14741 8960 14775
rect 8994 14741 9028 14775
rect 9062 14741 9096 14775
rect 9130 14741 9164 14775
rect 9198 14741 9232 14775
rect 9266 14741 9300 14775
rect 9334 14741 9368 14775
rect 9402 14741 9436 14775
rect 9470 14741 9504 14775
rect 9538 14741 9572 14775
rect 9606 14741 9640 14775
rect 9674 14741 9708 14775
rect 9742 14741 9776 14775
rect 9810 14741 9844 14775
rect 9878 14741 9912 14775
rect 9946 14741 9980 14775
rect 10014 14741 10048 14775
rect 10082 14741 10116 14775
rect 10150 14741 10184 14775
rect 10218 14741 10252 14775
rect 10286 14741 10320 14775
rect 10354 14741 10388 14775
rect 10422 14741 10456 14775
rect 10490 14741 10524 14775
rect 10558 14741 10592 14775
rect 10626 14741 10660 14775
rect 10694 14741 10728 14775
rect 10762 14741 10796 14775
rect 10830 14741 10864 14775
rect 10898 14741 10932 14775
rect 10966 14741 11000 14775
rect 11034 14741 11068 14775
rect 11102 14741 11136 14775
rect 11170 14741 11204 14775
rect 11238 14741 11272 14775
rect 11306 14741 11340 14775
rect 11374 14741 11408 14775
rect 11442 14741 11476 14775
rect 11510 14741 11544 14775
rect 11578 14741 11612 14775
rect 11646 14741 11680 14775
rect 11714 14741 11748 14775
rect 11782 14741 11816 14775
rect 11850 14741 11884 14775
rect 11918 14741 11952 14775
rect 11986 14741 12020 14775
rect 12054 14741 12088 14775
rect 12122 14741 12156 14775
rect 12190 14741 12224 14775
rect 12258 14741 12292 14775
rect 12326 14741 12360 14775
rect 12394 14741 12428 14775
rect 12462 14741 12496 14775
rect 12530 14741 12564 14775
rect 12598 14741 12632 14775
rect 12666 14741 12700 14775
rect 12734 14741 12768 14775
rect 12802 14741 12836 14775
rect 12870 14741 12904 14775
rect 12938 14741 12972 14775
rect 13006 14741 13040 14775
rect 13074 14741 13108 14775
rect 13142 14741 13176 14775
rect 13210 14741 13244 14775
rect 13278 14741 13312 14775
rect 13346 14741 13380 14775
rect 13414 14741 13448 14775
rect 13482 14741 13516 14775
rect 13550 14741 13584 14775
rect 13618 14741 13652 14775
rect 13686 14741 13720 14775
rect 13754 14741 13788 14775
rect 13822 14741 13856 14775
rect 13890 14741 13924 14775
rect 13958 14741 13992 14775
rect 14026 14741 14060 14775
rect 14094 14741 14128 14775
rect 14162 14741 14196 14775
<< locali >>
rect 245 36534 14724 36574
rect 245 36500 320 36534
rect 354 36533 14724 36534
rect 354 36500 14614 36533
rect 245 36499 14614 36500
rect 14648 36499 14724 36533
rect 245 36498 14724 36499
rect 245 36497 556 36498
rect 590 36497 628 36498
rect 662 36497 700 36498
rect 734 36497 772 36498
rect 806 36497 844 36498
rect 878 36497 916 36498
rect 950 36497 988 36498
rect 1022 36497 1060 36498
rect 1094 36497 1132 36498
rect 1166 36497 1204 36498
rect 1238 36497 1276 36498
rect 1310 36497 1348 36498
rect 1382 36497 1420 36498
rect 1454 36497 1492 36498
rect 1526 36497 1564 36498
rect 1598 36497 1636 36498
rect 1670 36497 1708 36498
rect 1742 36497 1780 36498
rect 1814 36497 1852 36498
rect 1886 36497 1924 36498
rect 1958 36497 1996 36498
rect 2030 36497 2068 36498
rect 2102 36497 2140 36498
rect 2174 36497 2212 36498
rect 2246 36497 2284 36498
rect 2318 36497 2356 36498
rect 2390 36497 2428 36498
rect 2462 36497 2500 36498
rect 2534 36497 2572 36498
rect 2606 36497 2644 36498
rect 2678 36497 2716 36498
rect 2750 36497 2788 36498
rect 2822 36497 2860 36498
rect 2894 36497 2932 36498
rect 2966 36497 3004 36498
rect 3038 36497 3076 36498
rect 3110 36497 3148 36498
rect 3182 36497 3220 36498
rect 3254 36497 3292 36498
rect 3326 36497 3364 36498
rect 3398 36497 3436 36498
rect 3470 36497 3508 36498
rect 3542 36497 3580 36498
rect 3614 36497 3652 36498
rect 3686 36497 3724 36498
rect 3758 36497 3796 36498
rect 3830 36497 3868 36498
rect 3902 36497 3940 36498
rect 3974 36497 4012 36498
rect 4046 36497 4084 36498
rect 4118 36497 4156 36498
rect 4190 36497 4228 36498
rect 4262 36497 4300 36498
rect 4334 36497 4372 36498
rect 4406 36497 4444 36498
rect 4478 36497 4516 36498
rect 4550 36497 4588 36498
rect 4622 36497 4660 36498
rect 4694 36497 4732 36498
rect 4766 36497 4804 36498
rect 4838 36497 4876 36498
rect 4910 36497 4948 36498
rect 4982 36497 5020 36498
rect 5054 36497 5092 36498
rect 5126 36497 5164 36498
rect 5198 36497 5236 36498
rect 5270 36497 5308 36498
rect 5342 36497 5380 36498
rect 5414 36497 5452 36498
rect 5486 36497 5524 36498
rect 5558 36497 5596 36498
rect 5630 36497 5668 36498
rect 5702 36497 5740 36498
rect 5774 36497 5812 36498
rect 5846 36497 5884 36498
rect 5918 36497 5956 36498
rect 5990 36497 6028 36498
rect 6062 36497 6100 36498
rect 6134 36497 6172 36498
rect 6206 36497 6244 36498
rect 6278 36497 6316 36498
rect 6350 36497 6388 36498
rect 6422 36497 6460 36498
rect 6494 36497 6532 36498
rect 6566 36497 6604 36498
rect 6638 36497 6676 36498
rect 6710 36497 6748 36498
rect 6782 36497 6820 36498
rect 6854 36497 6892 36498
rect 6926 36497 6964 36498
rect 6998 36497 7036 36498
rect 7070 36497 7108 36498
rect 7142 36497 7180 36498
rect 7214 36497 7252 36498
rect 7286 36497 7324 36498
rect 7358 36497 7396 36498
rect 7430 36497 7468 36498
rect 7502 36497 7540 36498
rect 7574 36497 7612 36498
rect 7646 36497 7684 36498
rect 7718 36497 7756 36498
rect 7790 36497 7828 36498
rect 7862 36497 7900 36498
rect 7934 36497 7972 36498
rect 8006 36497 8044 36498
rect 8078 36497 8116 36498
rect 8150 36497 8188 36498
rect 8222 36497 8260 36498
rect 8294 36497 8332 36498
rect 8366 36497 8404 36498
rect 8438 36497 8476 36498
rect 8510 36497 8548 36498
rect 8582 36497 8620 36498
rect 8654 36497 8692 36498
rect 8726 36497 8764 36498
rect 8798 36497 8836 36498
rect 8870 36497 8908 36498
rect 8942 36497 8980 36498
rect 9014 36497 9052 36498
rect 9086 36497 9124 36498
rect 9158 36497 9196 36498
rect 9230 36497 9268 36498
rect 9302 36497 9340 36498
rect 9374 36497 9412 36498
rect 9446 36497 9484 36498
rect 9518 36497 9556 36498
rect 9590 36497 9628 36498
rect 9662 36497 9700 36498
rect 9734 36497 9772 36498
rect 9806 36497 9844 36498
rect 9878 36497 9916 36498
rect 9950 36497 9988 36498
rect 10022 36497 10060 36498
rect 10094 36497 10132 36498
rect 10166 36497 10204 36498
rect 10238 36497 10276 36498
rect 10310 36497 10348 36498
rect 10382 36497 10420 36498
rect 10454 36497 10492 36498
rect 10526 36497 10564 36498
rect 10598 36497 10636 36498
rect 10670 36497 10708 36498
rect 10742 36497 10780 36498
rect 10814 36497 10852 36498
rect 10886 36497 10924 36498
rect 10958 36497 10996 36498
rect 11030 36497 11068 36498
rect 11102 36497 11140 36498
rect 11174 36497 11212 36498
rect 11246 36497 11284 36498
rect 11318 36497 11356 36498
rect 11390 36497 11428 36498
rect 11462 36497 11500 36498
rect 11534 36497 11572 36498
rect 11606 36497 11644 36498
rect 11678 36497 11716 36498
rect 11750 36497 11788 36498
rect 11822 36497 11860 36498
rect 11894 36497 11932 36498
rect 11966 36497 12004 36498
rect 12038 36497 12076 36498
rect 12110 36497 12148 36498
rect 12182 36497 12220 36498
rect 12254 36497 12292 36498
rect 12326 36497 12364 36498
rect 12398 36497 12436 36498
rect 12470 36497 12508 36498
rect 12542 36497 12580 36498
rect 12614 36497 12652 36498
rect 12686 36497 12724 36498
rect 12758 36497 12796 36498
rect 12830 36497 12868 36498
rect 12902 36497 12940 36498
rect 12974 36497 13012 36498
rect 13046 36497 13084 36498
rect 13118 36497 13156 36498
rect 13190 36497 13228 36498
rect 13262 36497 13300 36498
rect 13334 36497 13372 36498
rect 13406 36497 13444 36498
rect 13478 36497 13516 36498
rect 13550 36497 13588 36498
rect 13622 36497 13660 36498
rect 13694 36497 13732 36498
rect 13766 36497 13804 36498
rect 13838 36497 13876 36498
rect 13910 36497 13948 36498
rect 13982 36497 14020 36498
rect 14054 36497 14092 36498
rect 14126 36497 14164 36498
rect 14198 36497 14236 36498
rect 14270 36497 14308 36498
rect 14342 36497 14380 36498
rect 14414 36497 14724 36498
rect 245 36463 455 36497
rect 489 36463 523 36497
rect 590 36464 591 36497
rect 557 36463 591 36464
rect 625 36464 628 36497
rect 693 36464 700 36497
rect 761 36464 772 36497
rect 829 36464 844 36497
rect 897 36464 916 36497
rect 965 36464 988 36497
rect 1033 36464 1060 36497
rect 1101 36464 1132 36497
rect 625 36463 659 36464
rect 693 36463 727 36464
rect 761 36463 795 36464
rect 829 36463 863 36464
rect 897 36463 931 36464
rect 965 36463 999 36464
rect 1033 36463 1067 36464
rect 1101 36463 1135 36464
rect 1169 36463 1203 36497
rect 1238 36464 1271 36497
rect 1310 36464 1339 36497
rect 1382 36464 1407 36497
rect 1454 36464 1475 36497
rect 1526 36464 1543 36497
rect 1598 36464 1611 36497
rect 1670 36464 1679 36497
rect 1742 36464 1747 36497
rect 1814 36464 1815 36497
rect 1237 36463 1271 36464
rect 1305 36463 1339 36464
rect 1373 36463 1407 36464
rect 1441 36463 1475 36464
rect 1509 36463 1543 36464
rect 1577 36463 1611 36464
rect 1645 36463 1679 36464
rect 1713 36463 1747 36464
rect 1781 36463 1815 36464
rect 1849 36464 1852 36497
rect 1917 36464 1924 36497
rect 1985 36464 1996 36497
rect 2053 36464 2068 36497
rect 2121 36464 2140 36497
rect 2189 36464 2212 36497
rect 2257 36464 2284 36497
rect 2325 36464 2356 36497
rect 1849 36463 1883 36464
rect 1917 36463 1951 36464
rect 1985 36463 2019 36464
rect 2053 36463 2087 36464
rect 2121 36463 2155 36464
rect 2189 36463 2223 36464
rect 2257 36463 2291 36464
rect 2325 36463 2359 36464
rect 2393 36463 2427 36497
rect 2462 36464 2495 36497
rect 2534 36464 2563 36497
rect 2606 36464 2631 36497
rect 2678 36464 2699 36497
rect 2750 36464 2767 36497
rect 2822 36464 2835 36497
rect 2894 36464 2903 36497
rect 2966 36464 2971 36497
rect 3038 36464 3039 36497
rect 2461 36463 2495 36464
rect 2529 36463 2563 36464
rect 2597 36463 2631 36464
rect 2665 36463 2699 36464
rect 2733 36463 2767 36464
rect 2801 36463 2835 36464
rect 2869 36463 2903 36464
rect 2937 36463 2971 36464
rect 3005 36463 3039 36464
rect 3073 36464 3076 36497
rect 3141 36464 3148 36497
rect 3209 36464 3220 36497
rect 3277 36464 3292 36497
rect 3345 36464 3364 36497
rect 3413 36464 3436 36497
rect 3481 36464 3508 36497
rect 3549 36464 3580 36497
rect 3073 36463 3107 36464
rect 3141 36463 3175 36464
rect 3209 36463 3243 36464
rect 3277 36463 3311 36464
rect 3345 36463 3379 36464
rect 3413 36463 3447 36464
rect 3481 36463 3515 36464
rect 3549 36463 3583 36464
rect 3617 36463 3651 36497
rect 3686 36464 3719 36497
rect 3758 36464 3787 36497
rect 3830 36464 3855 36497
rect 3902 36464 3923 36497
rect 3974 36464 3991 36497
rect 4046 36464 4059 36497
rect 4118 36464 4127 36497
rect 4190 36464 4195 36497
rect 4262 36464 4263 36497
rect 3685 36463 3719 36464
rect 3753 36463 3787 36464
rect 3821 36463 3855 36464
rect 3889 36463 3923 36464
rect 3957 36463 3991 36464
rect 4025 36463 4059 36464
rect 4093 36463 4127 36464
rect 4161 36463 4195 36464
rect 4229 36463 4263 36464
rect 4297 36464 4300 36497
rect 4365 36464 4372 36497
rect 4433 36464 4444 36497
rect 4501 36464 4516 36497
rect 4569 36464 4588 36497
rect 4637 36464 4660 36497
rect 4705 36464 4732 36497
rect 4773 36464 4804 36497
rect 4297 36463 4331 36464
rect 4365 36463 4399 36464
rect 4433 36463 4467 36464
rect 4501 36463 4535 36464
rect 4569 36463 4603 36464
rect 4637 36463 4671 36464
rect 4705 36463 4739 36464
rect 4773 36463 4807 36464
rect 4841 36463 4875 36497
rect 4910 36464 4943 36497
rect 4982 36464 5011 36497
rect 5054 36464 5079 36497
rect 5126 36464 5147 36497
rect 5198 36464 5215 36497
rect 5270 36464 5283 36497
rect 5342 36464 5351 36497
rect 5414 36464 5419 36497
rect 5486 36464 5487 36497
rect 4909 36463 4943 36464
rect 4977 36463 5011 36464
rect 5045 36463 5079 36464
rect 5113 36463 5147 36464
rect 5181 36463 5215 36464
rect 5249 36463 5283 36464
rect 5317 36463 5351 36464
rect 5385 36463 5419 36464
rect 5453 36463 5487 36464
rect 5521 36464 5524 36497
rect 5589 36464 5596 36497
rect 5657 36464 5668 36497
rect 5725 36464 5740 36497
rect 5793 36464 5812 36497
rect 5861 36464 5884 36497
rect 5929 36464 5956 36497
rect 5997 36464 6028 36497
rect 5521 36463 5555 36464
rect 5589 36463 5623 36464
rect 5657 36463 5691 36464
rect 5725 36463 5759 36464
rect 5793 36463 5827 36464
rect 5861 36463 5895 36464
rect 5929 36463 5963 36464
rect 5997 36463 6031 36464
rect 6065 36463 6099 36497
rect 6134 36464 6167 36497
rect 6206 36464 6235 36497
rect 6278 36464 6303 36497
rect 6350 36464 6371 36497
rect 6422 36464 6439 36497
rect 6494 36464 6507 36497
rect 6566 36464 6575 36497
rect 6638 36464 6643 36497
rect 6710 36464 6711 36497
rect 6133 36463 6167 36464
rect 6201 36463 6235 36464
rect 6269 36463 6303 36464
rect 6337 36463 6371 36464
rect 6405 36463 6439 36464
rect 6473 36463 6507 36464
rect 6541 36463 6575 36464
rect 6609 36463 6643 36464
rect 6677 36463 6711 36464
rect 6745 36464 6748 36497
rect 6813 36464 6820 36497
rect 6881 36464 6892 36497
rect 6949 36464 6964 36497
rect 7017 36464 7036 36497
rect 7085 36464 7108 36497
rect 7153 36464 7180 36497
rect 7221 36464 7252 36497
rect 6745 36463 6779 36464
rect 6813 36463 6847 36464
rect 6881 36463 6915 36464
rect 6949 36463 6983 36464
rect 7017 36463 7051 36464
rect 7085 36463 7119 36464
rect 7153 36463 7187 36464
rect 7221 36463 7255 36464
rect 7289 36463 7323 36497
rect 7358 36464 7391 36497
rect 7430 36464 7459 36497
rect 7502 36464 7527 36497
rect 7574 36464 7595 36497
rect 7646 36464 7663 36497
rect 7718 36464 7731 36497
rect 7790 36464 7799 36497
rect 7862 36464 7867 36497
rect 7934 36464 7935 36497
rect 7357 36463 7391 36464
rect 7425 36463 7459 36464
rect 7493 36463 7527 36464
rect 7561 36463 7595 36464
rect 7629 36463 7663 36464
rect 7697 36463 7731 36464
rect 7765 36463 7799 36464
rect 7833 36463 7867 36464
rect 7901 36463 7935 36464
rect 7969 36464 7972 36497
rect 8037 36464 8044 36497
rect 8105 36464 8116 36497
rect 8173 36464 8188 36497
rect 8241 36464 8260 36497
rect 8309 36464 8332 36497
rect 8377 36464 8404 36497
rect 8445 36464 8476 36497
rect 7969 36463 8003 36464
rect 8037 36463 8071 36464
rect 8105 36463 8139 36464
rect 8173 36463 8207 36464
rect 8241 36463 8275 36464
rect 8309 36463 8343 36464
rect 8377 36463 8411 36464
rect 8445 36463 8479 36464
rect 8513 36463 8547 36497
rect 8582 36464 8615 36497
rect 8654 36464 8683 36497
rect 8726 36464 8751 36497
rect 8798 36464 8819 36497
rect 8870 36464 8887 36497
rect 8942 36464 8955 36497
rect 9014 36464 9023 36497
rect 9086 36464 9091 36497
rect 9158 36464 9159 36497
rect 8581 36463 8615 36464
rect 8649 36463 8683 36464
rect 8717 36463 8751 36464
rect 8785 36463 8819 36464
rect 8853 36463 8887 36464
rect 8921 36463 8955 36464
rect 8989 36463 9023 36464
rect 9057 36463 9091 36464
rect 9125 36463 9159 36464
rect 9193 36464 9196 36497
rect 9261 36464 9268 36497
rect 9329 36464 9340 36497
rect 9397 36464 9412 36497
rect 9465 36464 9484 36497
rect 9533 36464 9556 36497
rect 9601 36464 9628 36497
rect 9669 36464 9700 36497
rect 9193 36463 9227 36464
rect 9261 36463 9295 36464
rect 9329 36463 9363 36464
rect 9397 36463 9431 36464
rect 9465 36463 9499 36464
rect 9533 36463 9567 36464
rect 9601 36463 9635 36464
rect 9669 36463 9703 36464
rect 9737 36463 9771 36497
rect 9806 36464 9839 36497
rect 9878 36464 9907 36497
rect 9950 36464 9975 36497
rect 10022 36464 10043 36497
rect 10094 36464 10111 36497
rect 10166 36464 10179 36497
rect 10238 36464 10247 36497
rect 10310 36464 10315 36497
rect 10382 36464 10383 36497
rect 9805 36463 9839 36464
rect 9873 36463 9907 36464
rect 9941 36463 9975 36464
rect 10009 36463 10043 36464
rect 10077 36463 10111 36464
rect 10145 36463 10179 36464
rect 10213 36463 10247 36464
rect 10281 36463 10315 36464
rect 10349 36463 10383 36464
rect 10417 36464 10420 36497
rect 10485 36464 10492 36497
rect 10553 36464 10564 36497
rect 10621 36464 10636 36497
rect 10689 36464 10708 36497
rect 10757 36464 10780 36497
rect 10825 36464 10852 36497
rect 10893 36464 10924 36497
rect 10417 36463 10451 36464
rect 10485 36463 10519 36464
rect 10553 36463 10587 36464
rect 10621 36463 10655 36464
rect 10689 36463 10723 36464
rect 10757 36463 10791 36464
rect 10825 36463 10859 36464
rect 10893 36463 10927 36464
rect 10961 36463 10995 36497
rect 11030 36464 11063 36497
rect 11102 36464 11131 36497
rect 11174 36464 11199 36497
rect 11246 36464 11267 36497
rect 11318 36464 11335 36497
rect 11390 36464 11403 36497
rect 11462 36464 11471 36497
rect 11534 36464 11539 36497
rect 11606 36464 11607 36497
rect 11029 36463 11063 36464
rect 11097 36463 11131 36464
rect 11165 36463 11199 36464
rect 11233 36463 11267 36464
rect 11301 36463 11335 36464
rect 11369 36463 11403 36464
rect 11437 36463 11471 36464
rect 11505 36463 11539 36464
rect 11573 36463 11607 36464
rect 11641 36464 11644 36497
rect 11709 36464 11716 36497
rect 11777 36464 11788 36497
rect 11845 36464 11860 36497
rect 11913 36464 11932 36497
rect 11981 36464 12004 36497
rect 12049 36464 12076 36497
rect 12117 36464 12148 36497
rect 11641 36463 11675 36464
rect 11709 36463 11743 36464
rect 11777 36463 11811 36464
rect 11845 36463 11879 36464
rect 11913 36463 11947 36464
rect 11981 36463 12015 36464
rect 12049 36463 12083 36464
rect 12117 36463 12151 36464
rect 12185 36463 12219 36497
rect 12254 36464 12287 36497
rect 12326 36464 12355 36497
rect 12398 36464 12423 36497
rect 12470 36464 12491 36497
rect 12542 36464 12559 36497
rect 12614 36464 12627 36497
rect 12686 36464 12695 36497
rect 12758 36464 12763 36497
rect 12830 36464 12831 36497
rect 12253 36463 12287 36464
rect 12321 36463 12355 36464
rect 12389 36463 12423 36464
rect 12457 36463 12491 36464
rect 12525 36463 12559 36464
rect 12593 36463 12627 36464
rect 12661 36463 12695 36464
rect 12729 36463 12763 36464
rect 12797 36463 12831 36464
rect 12865 36464 12868 36497
rect 12933 36464 12940 36497
rect 13001 36464 13012 36497
rect 13069 36464 13084 36497
rect 13137 36464 13156 36497
rect 13205 36464 13228 36497
rect 13273 36464 13300 36497
rect 13341 36464 13372 36497
rect 12865 36463 12899 36464
rect 12933 36463 12967 36464
rect 13001 36463 13035 36464
rect 13069 36463 13103 36464
rect 13137 36463 13171 36464
rect 13205 36463 13239 36464
rect 13273 36463 13307 36464
rect 13341 36463 13375 36464
rect 13409 36463 13443 36497
rect 13478 36464 13511 36497
rect 13550 36464 13579 36497
rect 13622 36464 13647 36497
rect 13694 36464 13715 36497
rect 13766 36464 13783 36497
rect 13838 36464 13851 36497
rect 13910 36464 13919 36497
rect 13982 36464 13987 36497
rect 14054 36464 14055 36497
rect 13477 36463 13511 36464
rect 13545 36463 13579 36464
rect 13613 36463 13647 36464
rect 13681 36463 13715 36464
rect 13749 36463 13783 36464
rect 13817 36463 13851 36464
rect 13885 36463 13919 36464
rect 13953 36463 13987 36464
rect 14021 36463 14055 36464
rect 14089 36464 14092 36497
rect 14157 36464 14164 36497
rect 14225 36464 14236 36497
rect 14293 36464 14308 36497
rect 14361 36464 14380 36497
rect 14089 36463 14123 36464
rect 14157 36463 14191 36464
rect 14225 36463 14259 36464
rect 14293 36463 14327 36464
rect 14361 36463 14395 36464
rect 14429 36463 14463 36497
rect 14497 36463 14724 36497
rect 245 36462 14724 36463
rect 245 36428 320 36462
rect 354 36461 14724 36462
rect 354 36428 14614 36461
rect 245 36427 14614 36428
rect 14648 36427 14724 36461
rect 245 36389 14724 36427
rect 245 36356 430 36389
rect 245 36322 312 36356
rect 346 36322 430 36356
rect 245 36288 430 36322
rect 245 36254 312 36288
rect 346 36281 430 36288
rect 245 36247 320 36254
rect 354 36247 430 36281
rect 245 36220 430 36247
rect 245 36186 312 36220
rect 346 36209 430 36220
rect 245 36175 320 36186
rect 354 36175 430 36209
rect 14539 36362 14724 36389
rect 14539 36328 14607 36362
rect 14641 36328 14724 36362
rect 14539 36294 14724 36328
rect 14539 36260 14607 36294
rect 14641 36278 14724 36294
rect 14539 36244 14614 36260
rect 14648 36244 14724 36278
rect 14539 36226 14724 36244
rect 245 36152 430 36175
rect 245 36118 312 36152
rect 346 36137 430 36152
rect 245 36103 320 36118
rect 354 36103 430 36137
rect 245 36084 430 36103
rect 245 36050 312 36084
rect 346 36065 430 36084
rect 245 36031 320 36050
rect 354 36031 430 36065
rect 245 36016 430 36031
rect 245 35982 312 36016
rect 346 35993 430 36016
rect 245 35959 320 35982
rect 354 35959 430 35993
rect 245 35948 430 35959
rect 245 35914 312 35948
rect 346 35921 430 35948
rect 245 35887 320 35914
rect 354 35887 430 35921
rect 245 35880 430 35887
rect 245 35846 312 35880
rect 346 35849 430 35880
rect 245 35815 320 35846
rect 354 35815 430 35849
rect 245 35812 430 35815
rect 245 35778 312 35812
rect 346 35778 430 35812
rect 245 35777 430 35778
rect 245 35744 320 35777
rect 245 35710 312 35744
rect 354 35743 430 35777
rect 346 35710 430 35743
rect 245 35705 430 35710
rect 245 35676 320 35705
rect 245 35642 312 35676
rect 354 35671 430 35705
rect 346 35642 430 35671
rect 245 35633 430 35642
rect 245 35608 320 35633
rect 245 35574 312 35608
rect 354 35599 430 35633
rect 346 35574 430 35599
rect 245 35561 430 35574
rect 245 35540 320 35561
rect 245 35506 312 35540
rect 354 35527 430 35561
rect 346 35506 430 35527
rect 245 35489 430 35506
rect 245 35472 320 35489
rect 245 35438 312 35472
rect 354 35455 430 35489
rect 346 35438 430 35455
rect 245 35417 430 35438
rect 245 35404 320 35417
rect 245 35370 312 35404
rect 354 35383 430 35417
rect 346 35370 430 35383
rect 245 35345 430 35370
rect 245 35336 320 35345
rect 245 35302 312 35336
rect 354 35311 430 35345
rect 346 35302 430 35311
rect 245 35273 430 35302
rect 245 35268 320 35273
rect 245 35234 312 35268
rect 354 35239 430 35273
rect 346 35234 430 35239
rect 245 35201 430 35234
rect 245 35200 320 35201
rect 245 35166 312 35200
rect 354 35167 430 35201
rect 346 35166 430 35167
rect 245 35132 430 35166
rect 245 35098 312 35132
rect 346 35129 430 35132
rect 245 35095 320 35098
rect 354 35095 430 35129
rect 245 35064 430 35095
rect 245 35030 312 35064
rect 346 35057 430 35064
rect 245 35023 320 35030
rect 354 35023 430 35057
rect 245 34996 430 35023
rect 245 34962 312 34996
rect 346 34985 430 34996
rect 245 34951 320 34962
rect 354 34951 430 34985
rect 245 34928 430 34951
rect 245 34894 312 34928
rect 346 34913 430 34928
rect 245 34879 320 34894
rect 354 34879 430 34913
rect 245 34860 430 34879
rect 245 34826 312 34860
rect 346 34841 430 34860
rect 245 34807 320 34826
rect 354 34807 430 34841
rect 245 34792 430 34807
rect 245 34758 312 34792
rect 346 34769 430 34792
rect 245 34735 320 34758
rect 354 34735 430 34769
rect 245 34724 430 34735
rect 245 34690 312 34724
rect 346 34697 430 34724
rect 245 34663 320 34690
rect 354 34663 430 34697
rect 245 34656 430 34663
rect 245 34622 312 34656
rect 346 34625 430 34656
rect 245 34591 320 34622
rect 354 34591 430 34625
rect 245 34588 430 34591
rect 245 34554 312 34588
rect 346 34554 430 34588
rect 245 34553 430 34554
rect 245 34520 320 34553
rect 245 34486 312 34520
rect 354 34519 430 34553
rect 346 34486 430 34519
rect 245 34481 430 34486
rect 245 34452 320 34481
rect 245 34418 312 34452
rect 354 34447 430 34481
rect 346 34418 430 34447
rect 245 34409 430 34418
rect 245 34384 320 34409
rect 245 34350 312 34384
rect 354 34375 430 34409
rect 346 34350 430 34375
rect 245 34337 430 34350
rect 245 34316 320 34337
rect 245 34282 312 34316
rect 354 34303 430 34337
rect 346 34282 430 34303
rect 245 34265 430 34282
rect 245 34248 320 34265
rect 245 34214 312 34248
rect 354 34231 430 34265
rect 346 34214 430 34231
rect 245 34193 430 34214
rect 245 34180 320 34193
rect 245 34146 312 34180
rect 354 34159 430 34193
rect 346 34146 430 34159
rect 245 34121 430 34146
rect 245 34112 320 34121
rect 245 34078 312 34112
rect 354 34087 430 34121
rect 346 34078 430 34087
rect 245 34049 430 34078
rect 245 34044 320 34049
rect 245 34010 312 34044
rect 354 34015 430 34049
rect 346 34010 430 34015
rect 245 33977 430 34010
rect 245 33976 320 33977
rect 245 33942 312 33976
rect 354 33943 430 33977
rect 346 33942 430 33943
rect 245 33908 430 33942
rect 245 33874 312 33908
rect 346 33905 430 33908
rect 245 33871 320 33874
rect 354 33871 430 33905
rect 245 33840 430 33871
rect 245 33806 312 33840
rect 346 33833 430 33840
rect 245 33799 320 33806
rect 354 33799 430 33833
rect 245 33772 430 33799
rect 245 33738 312 33772
rect 346 33761 430 33772
rect 245 33727 320 33738
rect 354 33727 430 33761
rect 245 33704 430 33727
rect 245 33670 312 33704
rect 346 33689 430 33704
rect 245 33655 320 33670
rect 354 33655 430 33689
rect 245 33636 430 33655
rect 245 33602 312 33636
rect 346 33617 430 33636
rect 245 33583 320 33602
rect 354 33583 430 33617
rect 245 33568 430 33583
rect 245 33534 312 33568
rect 346 33545 430 33568
rect 245 33511 320 33534
rect 354 33511 430 33545
rect 245 33500 430 33511
rect 245 33466 312 33500
rect 346 33473 430 33500
rect 245 33439 320 33466
rect 354 33439 430 33473
rect 245 33432 430 33439
rect 245 33398 312 33432
rect 346 33401 430 33432
rect 245 33367 320 33398
rect 354 33367 430 33401
rect 245 33364 430 33367
rect 245 33330 312 33364
rect 346 33330 430 33364
rect 245 33329 430 33330
rect 245 33296 320 33329
rect 245 33262 312 33296
rect 354 33295 430 33329
rect 346 33262 430 33295
rect 245 33257 430 33262
rect 245 33228 320 33257
rect 245 33194 312 33228
rect 354 33223 430 33257
rect 346 33194 430 33223
rect 245 33185 430 33194
rect 245 33160 320 33185
rect 245 33126 312 33160
rect 354 33151 430 33185
rect 346 33126 430 33151
rect 245 33113 430 33126
rect 245 33092 320 33113
rect 245 33058 312 33092
rect 354 33079 430 33113
rect 346 33058 430 33079
rect 245 33041 430 33058
rect 245 33024 320 33041
rect 245 32990 312 33024
rect 354 33007 430 33041
rect 346 32990 430 33007
rect 245 32969 430 32990
rect 245 32956 320 32969
rect 245 32922 312 32956
rect 354 32935 430 32969
rect 346 32922 430 32935
rect 245 32897 430 32922
rect 245 32888 320 32897
rect 245 32854 312 32888
rect 354 32863 430 32897
rect 346 32854 430 32863
rect 245 32825 430 32854
rect 245 32820 320 32825
rect 245 32786 312 32820
rect 354 32791 430 32825
rect 346 32786 430 32791
rect 245 32753 430 32786
rect 245 32752 320 32753
rect 245 32718 312 32752
rect 354 32719 430 32753
rect 346 32718 430 32719
rect 245 32684 430 32718
rect 245 32650 312 32684
rect 346 32681 430 32684
rect 245 32647 320 32650
rect 354 32647 430 32681
rect 245 32616 430 32647
rect 245 32582 312 32616
rect 346 32609 430 32616
rect 245 32575 320 32582
rect 354 32575 430 32609
rect 245 32548 430 32575
rect 245 32514 312 32548
rect 346 32537 430 32548
rect 245 32503 320 32514
rect 354 32503 430 32537
rect 245 32480 430 32503
rect 245 32446 312 32480
rect 346 32465 430 32480
rect 245 32431 320 32446
rect 354 32431 430 32465
rect 245 32412 430 32431
rect 245 32378 312 32412
rect 346 32393 430 32412
rect 245 32359 320 32378
rect 354 32359 430 32393
rect 245 32344 430 32359
rect 245 32310 312 32344
rect 346 32321 430 32344
rect 245 32287 320 32310
rect 354 32287 430 32321
rect 245 32276 430 32287
rect 245 32242 312 32276
rect 346 32249 430 32276
rect 245 32215 320 32242
rect 354 32215 430 32249
rect 245 32208 430 32215
rect 245 32174 312 32208
rect 346 32177 430 32208
rect 245 32143 320 32174
rect 354 32143 430 32177
rect 245 32140 430 32143
rect 245 32106 312 32140
rect 346 32106 430 32140
rect 245 32105 430 32106
rect 245 32072 320 32105
rect 245 32038 312 32072
rect 354 32071 430 32105
rect 346 32038 430 32071
rect 245 32033 430 32038
rect 245 32004 320 32033
rect 245 31970 312 32004
rect 354 31999 430 32033
rect 346 31970 430 31999
rect 245 31961 430 31970
rect 245 31936 320 31961
rect 245 31902 312 31936
rect 354 31927 430 31961
rect 346 31902 430 31927
rect 245 31889 430 31902
rect 245 31868 320 31889
rect 245 31834 312 31868
rect 354 31855 430 31889
rect 346 31834 430 31855
rect 245 31817 430 31834
rect 245 31800 320 31817
rect 245 31766 312 31800
rect 354 31783 430 31817
rect 346 31766 430 31783
rect 245 31745 430 31766
rect 245 31732 320 31745
rect 245 31698 312 31732
rect 354 31711 430 31745
rect 346 31698 430 31711
rect 245 31673 430 31698
rect 245 31664 320 31673
rect 245 31630 312 31664
rect 354 31639 430 31673
rect 346 31630 430 31639
rect 245 31601 430 31630
rect 245 31596 320 31601
rect 245 31562 312 31596
rect 354 31567 430 31601
rect 346 31562 430 31567
rect 245 31529 430 31562
rect 245 31528 320 31529
rect 245 31494 312 31528
rect 354 31495 430 31529
rect 346 31494 430 31495
rect 245 31460 430 31494
rect 245 31426 312 31460
rect 346 31457 430 31460
rect 245 31423 320 31426
rect 354 31423 430 31457
rect 245 31392 430 31423
rect 245 31358 312 31392
rect 346 31385 430 31392
rect 245 31351 320 31358
rect 354 31351 430 31385
rect 245 31324 430 31351
rect 245 31290 312 31324
rect 346 31313 430 31324
rect 245 31279 320 31290
rect 354 31279 430 31313
rect 245 31256 430 31279
rect 245 31222 312 31256
rect 346 31241 430 31256
rect 245 31207 320 31222
rect 354 31207 430 31241
rect 245 31188 430 31207
rect 245 31154 312 31188
rect 346 31169 430 31188
rect 245 31135 320 31154
rect 354 31135 430 31169
rect 245 31120 430 31135
rect 245 31086 312 31120
rect 346 31097 430 31120
rect 245 31063 320 31086
rect 354 31063 430 31097
rect 245 31052 430 31063
rect 245 31018 312 31052
rect 346 31025 430 31052
rect 245 30991 320 31018
rect 354 30991 430 31025
rect 245 30984 430 30991
rect 245 30950 312 30984
rect 346 30953 430 30984
rect 245 30919 320 30950
rect 354 30919 430 30953
rect 245 30916 430 30919
rect 245 30882 312 30916
rect 346 30882 430 30916
rect 245 30881 430 30882
rect 245 30848 320 30881
rect 245 30814 312 30848
rect 354 30847 430 30881
rect 346 30814 430 30847
rect 245 30809 430 30814
rect 245 30780 320 30809
rect 245 30746 312 30780
rect 354 30775 430 30809
rect 346 30746 430 30775
rect 245 30737 430 30746
rect 245 30712 320 30737
rect 245 30678 312 30712
rect 354 30703 430 30737
rect 346 30678 430 30703
rect 245 30665 430 30678
rect 245 30644 320 30665
rect 245 30610 312 30644
rect 354 30631 430 30665
rect 346 30610 430 30631
rect 245 30593 430 30610
rect 245 30576 320 30593
rect 245 30542 312 30576
rect 354 30559 430 30593
rect 346 30542 430 30559
rect 245 30521 430 30542
rect 245 30508 320 30521
rect 245 30474 312 30508
rect 354 30487 430 30521
rect 346 30474 430 30487
rect 245 30449 430 30474
rect 245 30440 320 30449
rect 245 30406 312 30440
rect 354 30415 430 30449
rect 346 30406 430 30415
rect 245 30377 430 30406
rect 245 30372 320 30377
rect 245 30338 312 30372
rect 354 30343 430 30377
rect 346 30338 430 30343
rect 245 30305 430 30338
rect 245 30304 320 30305
rect 245 30270 312 30304
rect 354 30271 430 30305
rect 346 30270 430 30271
rect 245 30236 430 30270
rect 245 30202 312 30236
rect 346 30233 430 30236
rect 245 30199 320 30202
rect 354 30199 430 30233
rect 245 30168 430 30199
rect 245 30134 312 30168
rect 346 30161 430 30168
rect 245 30127 320 30134
rect 354 30127 430 30161
rect 245 30100 430 30127
rect 245 30066 312 30100
rect 346 30089 430 30100
rect 245 30055 320 30066
rect 354 30055 430 30089
rect 245 30032 430 30055
rect 245 29998 312 30032
rect 346 30017 430 30032
rect 245 29983 320 29998
rect 354 29983 430 30017
rect 245 29964 430 29983
rect 245 29930 312 29964
rect 346 29945 430 29964
rect 245 29911 320 29930
rect 354 29911 430 29945
rect 245 29896 430 29911
rect 245 29862 312 29896
rect 346 29873 430 29896
rect 245 29839 320 29862
rect 354 29839 430 29873
rect 245 29828 430 29839
rect 245 29794 312 29828
rect 346 29801 430 29828
rect 245 29767 320 29794
rect 354 29767 430 29801
rect 245 29760 430 29767
rect 245 29726 312 29760
rect 346 29729 430 29760
rect 245 29695 320 29726
rect 354 29695 430 29729
rect 245 29692 430 29695
rect 245 29658 312 29692
rect 346 29658 430 29692
rect 245 29657 430 29658
rect 245 29624 320 29657
rect 245 29590 312 29624
rect 354 29623 430 29657
rect 346 29590 430 29623
rect 245 29585 430 29590
rect 245 29556 320 29585
rect 245 29522 312 29556
rect 354 29551 430 29585
rect 346 29522 430 29551
rect 245 29513 430 29522
rect 245 29488 320 29513
rect 245 29454 312 29488
rect 354 29479 430 29513
rect 346 29454 430 29479
rect 245 29441 430 29454
rect 245 29420 320 29441
rect 245 29386 312 29420
rect 354 29407 430 29441
rect 346 29386 430 29407
rect 245 29369 430 29386
rect 245 29352 320 29369
rect 245 29318 312 29352
rect 354 29335 430 29369
rect 346 29318 430 29335
rect 245 29297 430 29318
rect 245 29284 320 29297
rect 245 29250 312 29284
rect 354 29263 430 29297
rect 346 29250 430 29263
rect 245 29225 430 29250
rect 245 29216 320 29225
rect 245 29182 312 29216
rect 354 29191 430 29225
rect 346 29182 430 29191
rect 245 29153 430 29182
rect 245 29148 320 29153
rect 245 29114 312 29148
rect 354 29119 430 29153
rect 346 29114 430 29119
rect 245 29081 430 29114
rect 245 29080 320 29081
rect 245 29046 312 29080
rect 354 29047 430 29081
rect 346 29046 430 29047
rect 245 29012 430 29046
rect 245 28978 312 29012
rect 346 29009 430 29012
rect 245 28975 320 28978
rect 354 28975 430 29009
rect 245 28944 430 28975
rect 245 28910 312 28944
rect 346 28937 430 28944
rect 245 28903 320 28910
rect 354 28903 430 28937
rect 245 28876 430 28903
rect 245 28842 312 28876
rect 346 28865 430 28876
rect 245 28831 320 28842
rect 354 28831 430 28865
rect 245 28808 430 28831
rect 245 28774 312 28808
rect 346 28793 430 28808
rect 245 28759 320 28774
rect 354 28759 430 28793
rect 245 28740 430 28759
rect 245 28706 312 28740
rect 346 28721 430 28740
rect 245 28687 320 28706
rect 354 28687 430 28721
rect 245 28672 430 28687
rect 245 28638 312 28672
rect 346 28649 430 28672
rect 245 28615 320 28638
rect 354 28615 430 28649
rect 245 28604 430 28615
rect 245 28570 312 28604
rect 346 28577 430 28604
rect 245 28543 320 28570
rect 354 28543 430 28577
rect 245 28536 430 28543
rect 245 28502 312 28536
rect 346 28505 430 28536
rect 245 28471 320 28502
rect 354 28471 430 28505
rect 245 28468 430 28471
rect 245 28434 312 28468
rect 346 28434 430 28468
rect 245 28433 430 28434
rect 245 28400 320 28433
rect 245 28366 312 28400
rect 354 28399 430 28433
rect 346 28366 430 28399
rect 245 28361 430 28366
rect 245 28332 320 28361
rect 245 28298 312 28332
rect 354 28327 430 28361
rect 346 28298 430 28327
rect 245 28289 430 28298
rect 245 28264 320 28289
rect 245 28230 312 28264
rect 354 28255 430 28289
rect 346 28230 430 28255
rect 245 28217 430 28230
rect 245 28196 320 28217
rect 245 28162 312 28196
rect 354 28183 430 28217
rect 346 28162 430 28183
rect 245 28145 430 28162
rect 245 28128 320 28145
rect 245 28094 312 28128
rect 354 28111 430 28145
rect 346 28094 430 28111
rect 245 28073 430 28094
rect 245 28060 320 28073
rect 245 28026 312 28060
rect 354 28039 430 28073
rect 346 28026 430 28039
rect 245 28001 430 28026
rect 245 27992 320 28001
rect 245 27958 312 27992
rect 354 27967 430 28001
rect 346 27958 430 27967
rect 245 27929 430 27958
rect 245 27924 320 27929
rect 245 27890 312 27924
rect 354 27895 430 27929
rect 346 27890 430 27895
rect 245 27857 430 27890
rect 245 27856 320 27857
rect 245 27822 312 27856
rect 354 27823 430 27857
rect 346 27822 430 27823
rect 245 27788 430 27822
rect 245 27754 312 27788
rect 346 27785 430 27788
rect 245 27751 320 27754
rect 354 27751 430 27785
rect 245 27720 430 27751
rect 245 27686 312 27720
rect 346 27713 430 27720
rect 245 27679 320 27686
rect 354 27679 430 27713
rect 245 27652 430 27679
rect 245 27618 312 27652
rect 346 27641 430 27652
rect 245 27607 320 27618
rect 354 27607 430 27641
rect 245 27584 430 27607
rect 245 27550 312 27584
rect 346 27569 430 27584
rect 245 27535 320 27550
rect 354 27535 430 27569
rect 245 27516 430 27535
rect 245 27482 312 27516
rect 346 27497 430 27516
rect 245 27463 320 27482
rect 354 27463 430 27497
rect 245 27448 430 27463
rect 245 27414 312 27448
rect 346 27425 430 27448
rect 245 27391 320 27414
rect 354 27391 430 27425
rect 245 27380 430 27391
rect 245 27346 312 27380
rect 346 27353 430 27380
rect 245 27319 320 27346
rect 354 27319 430 27353
rect 245 27312 430 27319
rect 245 27278 312 27312
rect 346 27281 430 27312
rect 245 27247 320 27278
rect 354 27247 430 27281
rect 245 27244 430 27247
rect 245 27210 312 27244
rect 346 27210 430 27244
rect 245 27209 430 27210
rect 245 27176 320 27209
rect 245 27142 312 27176
rect 354 27175 430 27209
rect 346 27142 430 27175
rect 245 27137 430 27142
rect 245 27108 320 27137
rect 245 27074 312 27108
rect 354 27103 430 27137
rect 346 27074 430 27103
rect 245 27065 430 27074
rect 245 27040 320 27065
rect 245 27006 312 27040
rect 354 27031 430 27065
rect 346 27006 430 27031
rect 245 26993 430 27006
rect 245 26972 320 26993
rect 245 26938 312 26972
rect 354 26959 430 26993
rect 346 26938 430 26959
rect 245 26921 430 26938
rect 245 26904 320 26921
rect 245 26870 312 26904
rect 354 26887 430 26921
rect 346 26870 430 26887
rect 245 26849 430 26870
rect 245 26836 320 26849
rect 245 26802 312 26836
rect 354 26815 430 26849
rect 346 26802 430 26815
rect 245 26777 430 26802
rect 245 26768 320 26777
rect 245 26734 312 26768
rect 354 26743 430 26777
rect 346 26734 430 26743
rect 245 26705 430 26734
rect 245 26700 320 26705
rect 245 26666 312 26700
rect 354 26671 430 26705
rect 346 26666 430 26671
rect 245 26633 430 26666
rect 245 26632 320 26633
rect 245 26598 312 26632
rect 354 26599 430 26633
rect 346 26598 430 26599
rect 245 26564 430 26598
rect 245 26530 312 26564
rect 346 26561 430 26564
rect 245 26527 320 26530
rect 354 26527 430 26561
rect 245 26496 430 26527
rect 245 26462 312 26496
rect 346 26489 430 26496
rect 245 26455 320 26462
rect 354 26455 430 26489
rect 245 26428 430 26455
rect 245 26394 312 26428
rect 346 26417 430 26428
rect 245 26383 320 26394
rect 354 26383 430 26417
rect 245 26360 430 26383
rect 245 26326 312 26360
rect 346 26345 430 26360
rect 245 26311 320 26326
rect 354 26311 430 26345
rect 245 26292 430 26311
rect 245 26258 312 26292
rect 346 26273 430 26292
rect 245 26239 320 26258
rect 354 26239 430 26273
rect 245 26224 430 26239
rect 245 26190 312 26224
rect 346 26201 430 26224
rect 245 26167 320 26190
rect 354 26167 430 26201
rect 245 26156 430 26167
rect 245 26122 312 26156
rect 346 26129 430 26156
rect 245 26095 320 26122
rect 354 26095 430 26129
rect 245 26088 430 26095
rect 245 26054 312 26088
rect 346 26057 430 26088
rect 245 26023 320 26054
rect 354 26023 430 26057
rect 245 26020 430 26023
rect 245 25986 312 26020
rect 346 25986 430 26020
rect 245 25985 430 25986
rect 245 25952 320 25985
rect 245 25918 312 25952
rect 354 25951 430 25985
rect 346 25918 430 25951
rect 245 25913 430 25918
rect 245 25884 320 25913
rect 245 25850 312 25884
rect 354 25879 430 25913
rect 346 25850 430 25879
rect 245 25841 430 25850
rect 245 25816 320 25841
rect 245 25782 312 25816
rect 354 25807 430 25841
rect 346 25782 430 25807
rect 245 25769 430 25782
rect 245 25748 320 25769
rect 245 25714 312 25748
rect 354 25735 430 25769
rect 346 25714 430 25735
rect 245 25697 430 25714
rect 245 25680 320 25697
rect 245 25646 312 25680
rect 354 25663 430 25697
rect 346 25646 430 25663
rect 245 25625 430 25646
rect 245 25612 320 25625
rect 245 25578 312 25612
rect 354 25591 430 25625
rect 346 25578 430 25591
rect 245 25553 430 25578
rect 245 25544 320 25553
rect 245 25510 312 25544
rect 354 25519 430 25553
rect 346 25510 430 25519
rect 245 25481 430 25510
rect 245 25476 320 25481
rect 245 25442 312 25476
rect 354 25447 430 25481
rect 346 25442 430 25447
rect 245 25409 430 25442
rect 245 25408 320 25409
rect 245 25374 312 25408
rect 354 25375 430 25409
rect 346 25374 430 25375
rect 245 25340 430 25374
rect 245 25306 312 25340
rect 346 25337 430 25340
rect 245 25303 320 25306
rect 354 25303 430 25337
rect 245 25272 430 25303
rect 245 25238 312 25272
rect 346 25265 430 25272
rect 245 25231 320 25238
rect 354 25231 430 25265
rect 245 25204 430 25231
rect 245 25170 312 25204
rect 346 25193 430 25204
rect 245 25159 320 25170
rect 354 25159 430 25193
rect 245 25136 430 25159
rect 245 25102 312 25136
rect 346 25121 430 25136
rect 245 25087 320 25102
rect 354 25087 430 25121
rect 245 25068 430 25087
rect 245 25034 312 25068
rect 346 25049 430 25068
rect 245 25015 320 25034
rect 354 25015 430 25049
rect 245 25000 430 25015
rect 245 24966 312 25000
rect 346 24977 430 25000
rect 245 24943 320 24966
rect 354 24943 430 24977
rect 245 24932 430 24943
rect 245 24898 312 24932
rect 346 24905 430 24932
rect 245 24871 320 24898
rect 354 24871 430 24905
rect 245 24864 430 24871
rect 245 24830 312 24864
rect 346 24833 430 24864
rect 245 24799 320 24830
rect 354 24799 430 24833
rect 245 24796 430 24799
rect 245 24762 312 24796
rect 346 24762 430 24796
rect 245 24761 430 24762
rect 245 24728 320 24761
rect 245 24694 312 24728
rect 354 24727 430 24761
rect 346 24694 430 24727
rect 245 24689 430 24694
rect 245 24660 320 24689
rect 245 24626 312 24660
rect 354 24655 430 24689
rect 346 24626 430 24655
rect 245 24617 430 24626
rect 245 24592 320 24617
rect 245 24558 312 24592
rect 354 24583 430 24617
rect 346 24558 430 24583
rect 245 24545 430 24558
rect 245 24524 320 24545
rect 245 24490 312 24524
rect 354 24511 430 24545
rect 346 24490 430 24511
rect 245 24473 430 24490
rect 245 24456 320 24473
rect 245 24422 312 24456
rect 354 24439 430 24473
rect 346 24422 430 24439
rect 245 24401 430 24422
rect 245 24388 320 24401
rect 245 24354 312 24388
rect 354 24367 430 24401
rect 346 24354 430 24367
rect 245 24329 430 24354
rect 245 24320 320 24329
rect 245 24286 312 24320
rect 354 24295 430 24329
rect 346 24286 430 24295
rect 245 24257 430 24286
rect 245 24252 320 24257
rect 245 24218 312 24252
rect 354 24223 430 24257
rect 346 24218 430 24223
rect 245 24185 430 24218
rect 245 24184 320 24185
rect 245 24150 312 24184
rect 354 24151 430 24185
rect 346 24150 430 24151
rect 245 24116 430 24150
rect 245 24082 312 24116
rect 346 24113 430 24116
rect 245 24079 320 24082
rect 354 24079 430 24113
rect 245 24048 430 24079
rect 245 24014 312 24048
rect 346 24041 430 24048
rect 245 24007 320 24014
rect 354 24007 430 24041
rect 245 23980 430 24007
rect 245 23946 312 23980
rect 346 23969 430 23980
rect 245 23935 320 23946
rect 354 23935 430 23969
rect 245 23912 430 23935
rect 245 23878 312 23912
rect 346 23897 430 23912
rect 245 23863 320 23878
rect 354 23863 430 23897
rect 245 23844 430 23863
rect 245 23810 312 23844
rect 346 23825 430 23844
rect 245 23791 320 23810
rect 354 23791 430 23825
rect 245 23776 430 23791
rect 245 23742 312 23776
rect 346 23753 430 23776
rect 245 23719 320 23742
rect 354 23719 430 23753
rect 245 23708 430 23719
rect 245 23674 312 23708
rect 346 23681 430 23708
rect 245 23647 320 23674
rect 354 23647 430 23681
rect 245 23640 430 23647
rect 245 23606 312 23640
rect 346 23609 430 23640
rect 245 23575 320 23606
rect 354 23575 430 23609
rect 245 23572 430 23575
rect 245 23538 312 23572
rect 346 23538 430 23572
rect 245 23537 430 23538
rect 245 23504 320 23537
rect 245 23470 312 23504
rect 354 23503 430 23537
rect 346 23470 430 23503
rect 245 23465 430 23470
rect 245 23436 320 23465
rect 245 23402 312 23436
rect 354 23431 430 23465
rect 346 23402 430 23431
rect 245 23393 430 23402
rect 245 23368 320 23393
rect 245 23334 312 23368
rect 354 23359 430 23393
rect 346 23334 430 23359
rect 245 23321 430 23334
rect 245 23300 320 23321
rect 245 23266 312 23300
rect 354 23287 430 23321
rect 346 23266 430 23287
rect 245 23249 430 23266
rect 245 23232 320 23249
rect 245 23198 312 23232
rect 354 23215 430 23249
rect 346 23198 430 23215
rect 245 23177 430 23198
rect 245 23164 320 23177
rect 245 23130 312 23164
rect 354 23143 430 23177
rect 346 23130 430 23143
rect 245 23105 430 23130
rect 245 23096 320 23105
rect 245 23062 312 23096
rect 354 23071 430 23105
rect 346 23062 430 23071
rect 245 23033 430 23062
rect 245 23028 320 23033
rect 245 22994 312 23028
rect 354 22999 430 23033
rect 346 22994 430 22999
rect 245 22961 430 22994
rect 245 22960 320 22961
rect 245 22926 312 22960
rect 354 22927 430 22961
rect 346 22926 430 22927
rect 245 22892 430 22926
rect 245 22858 312 22892
rect 346 22889 430 22892
rect 245 22855 320 22858
rect 354 22855 430 22889
rect 245 22824 430 22855
rect 245 22790 312 22824
rect 346 22817 430 22824
rect 245 22783 320 22790
rect 354 22783 430 22817
rect 245 22756 430 22783
rect 245 22722 312 22756
rect 346 22745 430 22756
rect 245 22711 320 22722
rect 354 22711 430 22745
rect 245 22688 430 22711
rect 245 22654 312 22688
rect 346 22673 430 22688
rect 245 22639 320 22654
rect 354 22639 430 22673
rect 245 22620 430 22639
rect 245 22586 312 22620
rect 346 22601 430 22620
rect 245 22567 320 22586
rect 354 22567 430 22601
rect 245 22552 430 22567
rect 245 22518 312 22552
rect 346 22529 430 22552
rect 245 22495 320 22518
rect 354 22495 430 22529
rect 245 22484 430 22495
rect 245 22450 312 22484
rect 346 22457 430 22484
rect 245 22423 320 22450
rect 354 22423 430 22457
rect 245 22416 430 22423
rect 245 22382 312 22416
rect 346 22385 430 22416
rect 245 22351 320 22382
rect 354 22351 430 22385
rect 245 22348 430 22351
rect 245 22314 312 22348
rect 346 22314 430 22348
rect 245 22313 430 22314
rect 245 22280 320 22313
rect 245 22246 312 22280
rect 354 22279 430 22313
rect 346 22246 430 22279
rect 245 22241 430 22246
rect 245 22212 320 22241
rect 245 22178 312 22212
rect 354 22207 430 22241
rect 346 22178 430 22207
rect 245 22169 430 22178
rect 245 22144 320 22169
rect 245 22110 312 22144
rect 354 22135 430 22169
rect 346 22110 430 22135
rect 245 22097 430 22110
rect 245 22076 320 22097
rect 245 22042 312 22076
rect 354 22063 430 22097
rect 346 22042 430 22063
rect 245 22025 430 22042
rect 245 22008 320 22025
rect 245 21974 312 22008
rect 354 21991 430 22025
rect 346 21974 430 21991
rect 245 21953 430 21974
rect 245 21940 320 21953
rect 245 21906 312 21940
rect 354 21919 430 21953
rect 346 21906 430 21919
rect 245 21881 430 21906
rect 245 21872 320 21881
rect 245 21838 312 21872
rect 354 21847 430 21881
rect 346 21838 430 21847
rect 245 21809 430 21838
rect 245 21804 320 21809
rect 245 21770 312 21804
rect 354 21775 430 21809
rect 346 21770 430 21775
rect 245 21737 430 21770
rect 245 21736 320 21737
rect 245 21702 312 21736
rect 354 21703 430 21737
rect 346 21702 430 21703
rect 245 21668 430 21702
rect 245 21634 312 21668
rect 346 21665 430 21668
rect 245 21631 320 21634
rect 354 21631 430 21665
rect 245 21600 430 21631
rect 245 21566 312 21600
rect 346 21593 430 21600
rect 245 21559 320 21566
rect 354 21559 430 21593
rect 245 21532 430 21559
rect 245 21498 312 21532
rect 346 21521 430 21532
rect 245 21487 320 21498
rect 354 21487 430 21521
rect 245 21464 430 21487
rect 245 21430 312 21464
rect 346 21449 430 21464
rect 245 21415 320 21430
rect 354 21415 430 21449
rect 245 21396 430 21415
rect 245 21362 312 21396
rect 346 21377 430 21396
rect 245 21343 320 21362
rect 354 21343 430 21377
rect 245 21328 430 21343
rect 245 21294 312 21328
rect 346 21305 430 21328
rect 245 21271 320 21294
rect 354 21271 430 21305
rect 245 21260 430 21271
rect 245 21226 312 21260
rect 346 21233 430 21260
rect 245 21199 320 21226
rect 354 21199 430 21233
rect 245 21192 430 21199
rect 245 21158 312 21192
rect 346 21161 430 21192
rect 245 21127 320 21158
rect 354 21127 430 21161
rect 245 21124 430 21127
rect 245 21090 312 21124
rect 346 21090 430 21124
rect 245 21089 430 21090
rect 245 21056 320 21089
rect 245 21022 312 21056
rect 354 21055 430 21089
rect 346 21022 430 21055
rect 245 21017 430 21022
rect 245 20988 320 21017
rect 245 20954 312 20988
rect 354 20983 430 21017
rect 346 20954 430 20983
rect 245 20945 430 20954
rect 245 20920 320 20945
rect 245 20886 312 20920
rect 354 20911 430 20945
rect 346 20886 430 20911
rect 245 20873 430 20886
rect 245 20852 320 20873
rect 245 20818 312 20852
rect 354 20839 430 20873
rect 346 20818 430 20839
rect 245 20801 430 20818
rect 245 20784 320 20801
rect 245 20750 312 20784
rect 354 20767 430 20801
rect 346 20750 430 20767
rect 245 20729 430 20750
rect 245 20716 320 20729
rect 245 20682 312 20716
rect 354 20695 430 20729
rect 346 20682 430 20695
rect 245 20657 430 20682
rect 245 20648 320 20657
rect 245 20614 312 20648
rect 354 20623 430 20657
rect 346 20614 430 20623
rect 245 20585 430 20614
rect 245 20580 320 20585
rect 245 20546 312 20580
rect 354 20551 430 20585
rect 346 20546 430 20551
rect 245 20513 430 20546
rect 245 20512 320 20513
rect 245 20478 312 20512
rect 354 20479 430 20513
rect 346 20478 430 20479
rect 245 20444 430 20478
rect 245 20410 312 20444
rect 346 20441 430 20444
rect 245 20407 320 20410
rect 354 20407 430 20441
rect 245 20376 430 20407
rect 245 20342 312 20376
rect 346 20369 430 20376
rect 245 20335 320 20342
rect 354 20335 430 20369
rect 245 20308 430 20335
rect 245 20274 312 20308
rect 346 20297 430 20308
rect 245 20263 320 20274
rect 354 20263 430 20297
rect 245 20240 430 20263
rect 245 20206 312 20240
rect 346 20225 430 20240
rect 245 20191 320 20206
rect 354 20191 430 20225
rect 245 20172 430 20191
rect 245 20138 312 20172
rect 346 20153 430 20172
rect 245 20119 320 20138
rect 354 20119 430 20153
rect 245 20104 430 20119
rect 245 20070 312 20104
rect 346 20081 430 20104
rect 245 20047 320 20070
rect 354 20047 430 20081
rect 245 20036 430 20047
rect 245 20002 312 20036
rect 346 20009 430 20036
rect 245 19975 320 20002
rect 354 19975 430 20009
rect 245 19968 430 19975
rect 245 19934 312 19968
rect 346 19937 430 19968
rect 245 19903 320 19934
rect 354 19903 430 19937
rect 245 19900 430 19903
rect 245 19866 312 19900
rect 346 19866 430 19900
rect 245 19865 430 19866
rect 245 19832 320 19865
rect 245 19798 312 19832
rect 354 19831 430 19865
rect 346 19798 430 19831
rect 245 19793 430 19798
rect 245 19764 320 19793
rect 245 19730 312 19764
rect 354 19759 430 19793
rect 346 19730 430 19759
rect 245 19721 430 19730
rect 245 19696 320 19721
rect 245 19662 312 19696
rect 354 19687 430 19721
rect 346 19662 430 19687
rect 245 19649 430 19662
rect 245 19628 320 19649
rect 245 19594 312 19628
rect 354 19615 430 19649
rect 346 19594 430 19615
rect 245 19577 430 19594
rect 245 19560 320 19577
rect 245 19526 312 19560
rect 354 19543 430 19577
rect 346 19526 430 19543
rect 245 19505 430 19526
rect 245 19492 320 19505
rect 245 19458 312 19492
rect 354 19471 430 19505
rect 346 19458 430 19471
rect 245 19433 430 19458
rect 245 19424 320 19433
rect 245 19390 312 19424
rect 354 19399 430 19433
rect 346 19390 430 19399
rect 245 19361 430 19390
rect 245 19356 320 19361
rect 245 19322 312 19356
rect 354 19327 430 19361
rect 346 19322 430 19327
rect 245 19289 430 19322
rect 245 19288 320 19289
rect 245 19254 312 19288
rect 354 19255 430 19289
rect 346 19254 430 19255
rect 245 19220 430 19254
rect 245 19186 312 19220
rect 346 19217 430 19220
rect 245 19183 320 19186
rect 354 19183 430 19217
rect 245 19152 430 19183
rect 245 19118 312 19152
rect 346 19145 430 19152
rect 245 19111 320 19118
rect 354 19111 430 19145
rect 245 19084 430 19111
rect 245 19050 312 19084
rect 346 19073 430 19084
rect 245 19039 320 19050
rect 354 19039 430 19073
rect 245 19016 430 19039
rect 245 18982 312 19016
rect 346 19001 430 19016
rect 245 18967 320 18982
rect 354 18967 430 19001
rect 245 18948 430 18967
rect 245 18914 312 18948
rect 346 18929 430 18948
rect 245 18895 320 18914
rect 354 18895 430 18929
rect 245 18880 430 18895
rect 245 18846 312 18880
rect 346 18857 430 18880
rect 245 18823 320 18846
rect 354 18823 430 18857
rect 245 18812 430 18823
rect 245 18778 312 18812
rect 346 18785 430 18812
rect 245 18751 320 18778
rect 354 18751 430 18785
rect 245 18744 430 18751
rect 245 18710 312 18744
rect 346 18713 430 18744
rect 245 18679 320 18710
rect 354 18679 430 18713
rect 245 18676 430 18679
rect 245 18642 312 18676
rect 346 18642 430 18676
rect 245 18641 430 18642
rect 245 18608 320 18641
rect 245 18574 312 18608
rect 354 18607 430 18641
rect 346 18574 430 18607
rect 245 18569 430 18574
rect 245 18540 320 18569
rect 245 18506 312 18540
rect 354 18535 430 18569
rect 346 18506 430 18535
rect 245 18497 430 18506
rect 245 18472 320 18497
rect 245 18438 312 18472
rect 354 18463 430 18497
rect 346 18438 430 18463
rect 245 18425 430 18438
rect 245 18404 320 18425
rect 245 18370 312 18404
rect 354 18391 430 18425
rect 346 18370 430 18391
rect 245 18353 430 18370
rect 245 18336 320 18353
rect 245 18302 312 18336
rect 354 18319 430 18353
rect 346 18302 430 18319
rect 245 18281 430 18302
rect 245 18268 320 18281
rect 245 18234 312 18268
rect 354 18247 430 18281
rect 346 18234 430 18247
rect 245 18209 430 18234
rect 245 18200 320 18209
rect 245 18166 312 18200
rect 354 18175 430 18209
rect 346 18166 430 18175
rect 245 18137 430 18166
rect 245 18132 320 18137
rect 245 18098 312 18132
rect 354 18103 430 18137
rect 346 18098 430 18103
rect 245 18065 430 18098
rect 245 18064 320 18065
rect 245 18030 312 18064
rect 354 18031 430 18065
rect 346 18030 430 18031
rect 245 17996 430 18030
rect 245 17962 312 17996
rect 346 17993 430 17996
rect 245 17959 320 17962
rect 354 17959 430 17993
rect 245 17928 430 17959
rect 245 17894 312 17928
rect 346 17921 430 17928
rect 245 17887 320 17894
rect 354 17887 430 17921
rect 245 17860 430 17887
rect 245 17826 312 17860
rect 346 17849 430 17860
rect 245 17815 320 17826
rect 354 17815 430 17849
rect 245 17792 430 17815
rect 245 17758 312 17792
rect 346 17777 430 17792
rect 245 17743 320 17758
rect 354 17743 430 17777
rect 245 17724 430 17743
rect 245 17690 312 17724
rect 346 17705 430 17724
rect 245 17671 320 17690
rect 354 17671 430 17705
rect 245 17656 430 17671
rect 245 17622 312 17656
rect 346 17633 430 17656
rect 245 17599 320 17622
rect 354 17599 430 17633
rect 245 17588 430 17599
rect 245 17554 312 17588
rect 346 17561 430 17588
rect 245 17527 320 17554
rect 354 17527 430 17561
rect 245 17520 430 17527
rect 245 17486 312 17520
rect 346 17489 430 17520
rect 245 17455 320 17486
rect 354 17455 430 17489
rect 245 17452 430 17455
rect 245 17418 312 17452
rect 346 17418 430 17452
rect 245 17417 430 17418
rect 245 17384 320 17417
rect 245 17350 312 17384
rect 354 17383 430 17417
rect 346 17350 430 17383
rect 245 17345 430 17350
rect 245 17316 320 17345
rect 245 17282 312 17316
rect 354 17311 430 17345
rect 346 17282 430 17311
rect 245 17273 430 17282
rect 245 17248 320 17273
rect 245 17214 312 17248
rect 354 17239 430 17273
rect 346 17214 430 17239
rect 245 17201 430 17214
rect 245 17180 320 17201
rect 245 17146 312 17180
rect 354 17167 430 17201
rect 346 17146 430 17167
rect 245 17129 430 17146
rect 245 17112 320 17129
rect 245 17078 312 17112
rect 354 17095 430 17129
rect 346 17078 430 17095
rect 245 17057 430 17078
rect 245 17044 320 17057
rect 245 17010 312 17044
rect 354 17023 430 17057
rect 346 17010 430 17023
rect 245 16985 430 17010
rect 245 16976 320 16985
rect 245 16942 312 16976
rect 354 16951 430 16985
rect 346 16942 430 16951
rect 245 16913 430 16942
rect 245 16908 320 16913
rect 245 16874 312 16908
rect 354 16879 430 16913
rect 346 16874 430 16879
rect 245 16841 430 16874
rect 245 16840 320 16841
rect 245 16806 312 16840
rect 354 16807 430 16841
rect 346 16806 430 16807
rect 245 16772 430 16806
rect 245 16738 312 16772
rect 346 16769 430 16772
rect 245 16735 320 16738
rect 354 16735 430 16769
rect 245 16704 430 16735
rect 245 16670 312 16704
rect 346 16697 430 16704
rect 245 16663 320 16670
rect 354 16663 430 16697
rect 245 16636 430 16663
rect 245 16602 312 16636
rect 346 16625 430 16636
rect 245 16591 320 16602
rect 354 16591 430 16625
rect 245 16568 430 16591
rect 245 16534 312 16568
rect 346 16553 430 16568
rect 245 16519 320 16534
rect 354 16519 430 16553
rect 245 16500 430 16519
rect 245 16466 312 16500
rect 346 16481 430 16500
rect 245 16447 320 16466
rect 354 16447 430 16481
rect 245 16432 430 16447
rect 245 16398 312 16432
rect 346 16409 430 16432
rect 245 16375 320 16398
rect 354 16375 430 16409
rect 245 16364 430 16375
rect 245 16330 312 16364
rect 346 16337 430 16364
rect 245 16303 320 16330
rect 354 16303 430 16337
rect 245 16296 430 16303
rect 245 16262 312 16296
rect 346 16265 430 16296
rect 245 16231 320 16262
rect 354 16231 430 16265
rect 245 16228 430 16231
rect 245 16194 312 16228
rect 346 16194 430 16228
rect 245 16193 430 16194
rect 245 16160 320 16193
rect 245 16126 312 16160
rect 354 16159 430 16193
rect 346 16126 430 16159
rect 245 16121 430 16126
rect 245 16092 320 16121
rect 245 16058 312 16092
rect 354 16087 430 16121
rect 346 16058 430 16087
rect 245 16049 430 16058
rect 245 16024 320 16049
rect 245 15990 312 16024
rect 354 16015 430 16049
rect 346 15990 430 16015
rect 245 15977 430 15990
rect 245 15956 320 15977
rect 245 15922 312 15956
rect 354 15943 430 15977
rect 346 15922 430 15943
rect 245 15905 430 15922
rect 245 15888 320 15905
rect 245 15854 312 15888
rect 354 15871 430 15905
rect 346 15854 430 15871
rect 245 15833 430 15854
rect 245 15820 320 15833
rect 245 15786 312 15820
rect 354 15799 430 15833
rect 346 15786 430 15799
rect 245 15761 430 15786
rect 245 15752 320 15761
rect 245 15718 312 15752
rect 354 15727 430 15761
rect 346 15718 430 15727
rect 245 15689 430 15718
rect 245 15684 320 15689
rect 245 15650 312 15684
rect 354 15655 430 15689
rect 346 15650 430 15655
rect 245 15617 430 15650
rect 245 15616 320 15617
rect 245 15582 312 15616
rect 354 15583 430 15617
rect 346 15582 430 15583
rect 245 15548 430 15582
rect 245 15514 312 15548
rect 346 15545 430 15548
rect 245 15511 320 15514
rect 354 15511 430 15545
rect 245 15480 430 15511
rect 245 15446 312 15480
rect 346 15473 430 15480
rect 245 15439 320 15446
rect 354 15439 430 15473
rect 245 15412 430 15439
rect 245 15378 312 15412
rect 346 15401 430 15412
rect 245 15367 320 15378
rect 354 15367 430 15401
rect 245 15344 430 15367
rect 245 15310 312 15344
rect 346 15329 430 15344
rect 245 15295 320 15310
rect 354 15295 430 15329
rect 245 15276 430 15295
rect 245 15242 312 15276
rect 346 15257 430 15276
rect 245 15223 320 15242
rect 354 15223 430 15257
rect 245 15208 430 15223
rect 245 15174 312 15208
rect 346 15185 430 15208
rect 245 15151 320 15174
rect 354 15151 430 15185
rect 245 15140 430 15151
rect 245 15106 312 15140
rect 346 15113 430 15140
rect 245 15079 320 15106
rect 354 15079 430 15113
rect 245 15072 430 15079
rect 245 15038 312 15072
rect 346 15041 430 15072
rect 245 15007 320 15038
rect 354 15007 430 15041
rect 245 15004 430 15007
rect 245 14970 312 15004
rect 346 14970 430 15004
rect 245 14969 430 14970
rect 245 14936 320 14969
rect 245 14902 312 14936
rect 354 14935 430 14969
rect 346 14902 430 14935
rect 245 14897 430 14902
rect 245 14868 320 14897
rect 245 14834 312 14868
rect 354 14863 430 14897
rect 346 14834 430 14863
rect 245 14825 430 14834
rect 245 14800 320 14825
rect 245 14766 312 14800
rect 354 14791 430 14825
rect 346 14766 430 14791
rect 245 14753 430 14766
rect 245 14732 320 14753
rect 245 14698 312 14732
rect 354 14719 430 14753
rect 346 14698 430 14719
rect 603 36177 14361 36207
rect 603 36143 766 36177
rect 800 36143 834 36177
rect 868 36143 902 36177
rect 936 36143 970 36177
rect 1004 36143 1038 36177
rect 1072 36143 1106 36177
rect 1140 36143 1174 36177
rect 1208 36143 1242 36177
rect 1276 36143 1310 36177
rect 1344 36143 1378 36177
rect 1412 36143 1446 36177
rect 1480 36143 1514 36177
rect 1548 36143 1582 36177
rect 1616 36143 1650 36177
rect 1684 36143 1718 36177
rect 1752 36143 1786 36177
rect 1820 36143 1854 36177
rect 1888 36143 1922 36177
rect 1956 36143 1990 36177
rect 2024 36143 2058 36177
rect 2092 36143 2126 36177
rect 2160 36143 2194 36177
rect 2228 36143 2262 36177
rect 2296 36143 2330 36177
rect 2364 36143 2398 36177
rect 2432 36143 2466 36177
rect 2500 36143 2534 36177
rect 2568 36143 2602 36177
rect 2636 36143 2670 36177
rect 2704 36143 2738 36177
rect 2772 36143 2806 36177
rect 2840 36143 2874 36177
rect 2908 36143 2942 36177
rect 2976 36143 3010 36177
rect 3044 36143 3078 36177
rect 3112 36143 3146 36177
rect 3180 36143 3214 36177
rect 3248 36143 3282 36177
rect 3316 36143 3350 36177
rect 3384 36143 3418 36177
rect 3452 36143 3486 36177
rect 3520 36143 3554 36177
rect 3588 36143 3622 36177
rect 3656 36143 3690 36177
rect 3724 36143 3758 36177
rect 3792 36143 3826 36177
rect 3860 36143 3894 36177
rect 3928 36143 3962 36177
rect 3996 36143 4030 36177
rect 4064 36143 4098 36177
rect 4132 36143 4166 36177
rect 4200 36143 4234 36177
rect 4268 36143 4302 36177
rect 4336 36143 4370 36177
rect 4404 36143 4438 36177
rect 4472 36143 4506 36177
rect 4540 36143 4574 36177
rect 4608 36143 4642 36177
rect 4676 36143 4710 36177
rect 4744 36143 4778 36177
rect 4812 36143 4846 36177
rect 4880 36143 4914 36177
rect 4948 36143 4982 36177
rect 5016 36143 5050 36177
rect 5084 36143 5118 36177
rect 5152 36143 5186 36177
rect 5220 36143 5254 36177
rect 5288 36143 5322 36177
rect 5356 36143 5390 36177
rect 5424 36143 5458 36177
rect 5492 36143 5526 36177
rect 5560 36143 5594 36177
rect 5628 36143 5662 36177
rect 5696 36143 5730 36177
rect 5764 36143 5798 36177
rect 5832 36143 5866 36177
rect 5900 36143 5934 36177
rect 5968 36143 6002 36177
rect 6036 36143 6070 36177
rect 6104 36143 6138 36177
rect 6172 36143 6206 36177
rect 6240 36143 6274 36177
rect 6308 36143 6342 36177
rect 6376 36143 6410 36177
rect 6444 36143 6478 36177
rect 6512 36143 6546 36177
rect 6580 36143 6614 36177
rect 6648 36143 6682 36177
rect 6716 36143 6750 36177
rect 6784 36143 6818 36177
rect 6852 36143 6886 36177
rect 6920 36143 6954 36177
rect 6988 36143 7022 36177
rect 7056 36143 7090 36177
rect 7124 36143 7158 36177
rect 7192 36143 7226 36177
rect 7260 36143 7294 36177
rect 7328 36143 7362 36177
rect 7396 36143 7430 36177
rect 7464 36143 7498 36177
rect 7532 36143 7566 36177
rect 7600 36143 7634 36177
rect 7668 36143 7702 36177
rect 7736 36143 7770 36177
rect 7804 36143 7838 36177
rect 7872 36143 7906 36177
rect 7940 36143 7974 36177
rect 8008 36143 8042 36177
rect 8076 36143 8110 36177
rect 8144 36143 8178 36177
rect 8212 36143 8246 36177
rect 8280 36143 8314 36177
rect 8348 36143 8382 36177
rect 8416 36143 8450 36177
rect 8484 36143 8518 36177
rect 8552 36143 8586 36177
rect 8620 36143 8654 36177
rect 8688 36143 8722 36177
rect 8756 36143 8790 36177
rect 8824 36143 8858 36177
rect 8892 36143 8926 36177
rect 8960 36143 8994 36177
rect 9028 36143 9062 36177
rect 9096 36143 9130 36177
rect 9164 36143 9198 36177
rect 9232 36143 9266 36177
rect 9300 36143 9334 36177
rect 9368 36143 9402 36177
rect 9436 36143 9470 36177
rect 9504 36143 9538 36177
rect 9572 36143 9606 36177
rect 9640 36143 9674 36177
rect 9708 36143 9742 36177
rect 9776 36143 9810 36177
rect 9844 36143 9878 36177
rect 9912 36143 9946 36177
rect 9980 36143 10014 36177
rect 10048 36143 10082 36177
rect 10116 36143 10150 36177
rect 10184 36143 10218 36177
rect 10252 36143 10286 36177
rect 10320 36143 10354 36177
rect 10388 36143 10422 36177
rect 10456 36143 10490 36177
rect 10524 36143 10558 36177
rect 10592 36143 10626 36177
rect 10660 36143 10694 36177
rect 10728 36143 10762 36177
rect 10796 36143 10830 36177
rect 10864 36143 10898 36177
rect 10932 36143 10966 36177
rect 11000 36143 11034 36177
rect 11068 36143 11102 36177
rect 11136 36143 11170 36177
rect 11204 36143 11238 36177
rect 11272 36143 11306 36177
rect 11340 36143 11374 36177
rect 11408 36143 11442 36177
rect 11476 36143 11510 36177
rect 11544 36143 11578 36177
rect 11612 36143 11646 36177
rect 11680 36143 11714 36177
rect 11748 36143 11782 36177
rect 11816 36143 11850 36177
rect 11884 36143 11918 36177
rect 11952 36143 11986 36177
rect 12020 36143 12054 36177
rect 12088 36143 12122 36177
rect 12156 36143 12190 36177
rect 12224 36143 12258 36177
rect 12292 36143 12326 36177
rect 12360 36143 12394 36177
rect 12428 36143 12462 36177
rect 12496 36143 12530 36177
rect 12564 36143 12598 36177
rect 12632 36143 12666 36177
rect 12700 36143 12734 36177
rect 12768 36143 12802 36177
rect 12836 36143 12870 36177
rect 12904 36143 12938 36177
rect 12972 36143 13006 36177
rect 13040 36143 13074 36177
rect 13108 36143 13142 36177
rect 13176 36143 13210 36177
rect 13244 36143 13278 36177
rect 13312 36143 13346 36177
rect 13380 36143 13414 36177
rect 13448 36143 13482 36177
rect 13516 36143 13550 36177
rect 13584 36143 13618 36177
rect 13652 36143 13686 36177
rect 13720 36143 13754 36177
rect 13788 36143 13822 36177
rect 13856 36143 13890 36177
rect 13924 36143 13958 36177
rect 13992 36143 14026 36177
rect 14060 36143 14094 36177
rect 14128 36143 14162 36177
rect 14196 36143 14361 36177
rect 603 36050 14361 36143
rect 603 36016 632 36050
rect 666 36016 14297 36050
rect 14331 36016 14361 36050
rect 603 36003 14361 36016
rect 603 35982 1009 36003
rect 603 35948 632 35982
rect 666 35969 1009 35982
rect 1043 35969 1081 36003
rect 1115 35969 1153 36003
rect 1187 35969 1225 36003
rect 1259 35969 1297 36003
rect 1331 35969 1369 36003
rect 1403 35969 1441 36003
rect 1475 35969 1513 36003
rect 1547 35969 1585 36003
rect 1619 35969 1657 36003
rect 1691 35969 1729 36003
rect 1763 35969 1801 36003
rect 1835 35969 1873 36003
rect 1907 35969 1945 36003
rect 1979 35969 2017 36003
rect 2051 35969 2089 36003
rect 2123 35969 2161 36003
rect 2195 35969 2233 36003
rect 2267 35969 2305 36003
rect 2339 35969 2377 36003
rect 2411 35969 2449 36003
rect 2483 35969 2521 36003
rect 2555 35969 2593 36003
rect 2627 35969 2665 36003
rect 2699 35969 2737 36003
rect 2771 35969 2809 36003
rect 2843 35969 2881 36003
rect 2915 35969 2953 36003
rect 2987 35969 3025 36003
rect 3059 35969 3097 36003
rect 3131 35969 3169 36003
rect 3203 35969 3241 36003
rect 3275 35969 3313 36003
rect 3347 35969 3385 36003
rect 3419 35969 3457 36003
rect 3491 35969 3529 36003
rect 3563 35969 3601 36003
rect 3635 35969 3673 36003
rect 3707 35969 3745 36003
rect 3779 35969 3817 36003
rect 3851 35969 3889 36003
rect 3923 35969 3961 36003
rect 3995 35969 4033 36003
rect 4067 35969 4105 36003
rect 4139 35969 4177 36003
rect 4211 35969 4249 36003
rect 4283 35969 4321 36003
rect 4355 35969 4393 36003
rect 4427 35969 4465 36003
rect 4499 35969 4537 36003
rect 4571 35969 4609 36003
rect 4643 35969 4681 36003
rect 4715 35969 4753 36003
rect 4787 35969 4825 36003
rect 4859 35969 4897 36003
rect 4931 35969 4969 36003
rect 5003 35969 5041 36003
rect 5075 35969 5113 36003
rect 5147 35969 5185 36003
rect 5219 35969 5257 36003
rect 5291 35969 5329 36003
rect 5363 35969 5401 36003
rect 5435 35969 5473 36003
rect 5507 35969 5545 36003
rect 5579 35969 5617 36003
rect 5651 35969 5689 36003
rect 5723 35969 5761 36003
rect 5795 35969 5833 36003
rect 5867 35969 5905 36003
rect 5939 35969 5977 36003
rect 6011 35969 6049 36003
rect 6083 35969 6121 36003
rect 6155 35969 6193 36003
rect 6227 35969 6265 36003
rect 6299 35969 6337 36003
rect 6371 35969 6409 36003
rect 6443 35969 6481 36003
rect 6515 35969 6553 36003
rect 6587 35969 6625 36003
rect 6659 35969 6697 36003
rect 6731 35969 6769 36003
rect 6803 35969 6841 36003
rect 6875 35969 6913 36003
rect 6947 35969 6985 36003
rect 7019 35969 7057 36003
rect 7091 35969 7129 36003
rect 7163 35969 7201 36003
rect 7235 35969 7273 36003
rect 7307 35969 7345 36003
rect 7379 35969 7417 36003
rect 7451 35969 7489 36003
rect 7523 35969 7561 36003
rect 7595 35969 7633 36003
rect 7667 35969 7705 36003
rect 7739 35969 7777 36003
rect 7811 35969 7849 36003
rect 7883 35969 7921 36003
rect 7955 35969 7993 36003
rect 8027 35969 8065 36003
rect 8099 35969 8137 36003
rect 8171 35969 8209 36003
rect 8243 35969 8281 36003
rect 8315 35969 8353 36003
rect 8387 35969 8425 36003
rect 8459 35969 8497 36003
rect 8531 35969 8569 36003
rect 8603 35969 8641 36003
rect 8675 35969 8713 36003
rect 8747 35969 8785 36003
rect 8819 35969 8857 36003
rect 8891 35969 8929 36003
rect 8963 35969 9001 36003
rect 9035 35969 9073 36003
rect 9107 35969 9145 36003
rect 9179 35969 9217 36003
rect 9251 35969 9289 36003
rect 9323 35969 9361 36003
rect 9395 35969 9433 36003
rect 9467 35969 9505 36003
rect 9539 35969 9577 36003
rect 9611 35969 9649 36003
rect 9683 35969 9721 36003
rect 9755 35969 9793 36003
rect 9827 35969 9865 36003
rect 9899 35969 9937 36003
rect 9971 35969 10009 36003
rect 10043 35969 10081 36003
rect 10115 35969 10153 36003
rect 10187 35969 10225 36003
rect 10259 35969 10297 36003
rect 10331 35969 10369 36003
rect 10403 35969 10441 36003
rect 10475 35969 10513 36003
rect 10547 35969 10585 36003
rect 10619 35969 10657 36003
rect 10691 35969 10729 36003
rect 10763 35969 10801 36003
rect 10835 35969 10873 36003
rect 10907 35969 10945 36003
rect 10979 35969 11017 36003
rect 11051 35969 11089 36003
rect 11123 35969 11161 36003
rect 11195 35969 11233 36003
rect 11267 35969 11305 36003
rect 11339 35969 11377 36003
rect 11411 35969 11449 36003
rect 11483 35969 11521 36003
rect 11555 35969 11593 36003
rect 11627 35969 11665 36003
rect 11699 35969 11737 36003
rect 11771 35969 11809 36003
rect 11843 35969 11881 36003
rect 11915 35969 11953 36003
rect 11987 35969 12025 36003
rect 12059 35969 12097 36003
rect 12131 35969 12169 36003
rect 12203 35969 12241 36003
rect 12275 35969 12313 36003
rect 12347 35969 12385 36003
rect 12419 35969 12457 36003
rect 12491 35969 12529 36003
rect 12563 35969 12601 36003
rect 12635 35969 12673 36003
rect 12707 35969 12745 36003
rect 12779 35969 12817 36003
rect 12851 35969 12889 36003
rect 12923 35969 12961 36003
rect 12995 35969 13033 36003
rect 13067 35969 13105 36003
rect 13139 35969 13177 36003
rect 13211 35969 13249 36003
rect 13283 35969 13321 36003
rect 13355 35969 13393 36003
rect 13427 35969 13465 36003
rect 13499 35969 13537 36003
rect 13571 35969 13609 36003
rect 13643 35969 13681 36003
rect 13715 35969 13753 36003
rect 13787 35969 13825 36003
rect 13859 35969 13897 36003
rect 13931 35969 13969 36003
rect 14003 35982 14361 36003
rect 14003 35969 14297 35982
rect 666 35948 14297 35969
rect 14331 35948 14361 35982
rect 603 35914 14361 35948
rect 603 35880 632 35914
rect 666 35900 14297 35914
rect 666 35880 807 35900
rect 603 35866 807 35880
rect 841 35880 14297 35900
rect 14331 35880 14361 35914
rect 841 35866 14361 35880
rect 603 35846 14361 35866
rect 603 35812 632 35846
rect 666 35828 14297 35846
rect 666 35812 807 35828
rect 603 35794 807 35812
rect 841 35821 14297 35828
rect 841 35794 14122 35821
rect 603 35787 14122 35794
rect 14156 35812 14297 35821
rect 14331 35812 14361 35846
rect 14156 35787 14361 35812
rect 603 35778 14361 35787
rect 603 35744 632 35778
rect 666 35756 14297 35778
rect 666 35744 807 35756
rect 603 35722 807 35744
rect 841 35749 14297 35756
rect 841 35722 14122 35749
rect 603 35715 14122 35722
rect 14156 35744 14297 35749
rect 14331 35744 14361 35778
rect 14156 35715 14361 35744
rect 603 35710 14361 35715
rect 603 35676 632 35710
rect 666 35684 14297 35710
rect 666 35676 807 35684
rect 603 35650 807 35676
rect 841 35677 14297 35684
rect 841 35650 14122 35677
rect 603 35643 14122 35650
rect 14156 35676 14297 35677
rect 14331 35676 14361 35710
rect 14156 35643 14361 35676
rect 603 35642 14361 35643
rect 603 35608 632 35642
rect 666 35612 14297 35642
rect 666 35608 807 35612
rect 603 35578 807 35608
rect 841 35608 14297 35612
rect 14331 35608 14361 35642
rect 841 35605 14361 35608
rect 841 35578 14122 35605
rect 603 35574 14122 35578
rect 603 35540 632 35574
rect 666 35571 14122 35574
rect 14156 35574 14361 35605
rect 14156 35571 14297 35574
rect 666 35540 14297 35571
rect 14331 35540 14361 35574
rect 603 35506 807 35540
rect 841 35533 14361 35540
rect 841 35506 14122 35533
rect 603 35472 632 35506
rect 666 35499 14122 35506
rect 14156 35506 14361 35533
rect 14156 35499 14297 35506
rect 666 35472 14297 35499
rect 14331 35472 14361 35506
rect 603 35468 14361 35472
rect 603 35438 807 35468
rect 603 35404 632 35438
rect 666 35434 807 35438
rect 841 35461 14361 35468
rect 841 35434 14122 35461
rect 666 35427 14122 35434
rect 14156 35438 14361 35461
rect 14156 35427 14297 35438
rect 666 35404 14297 35427
rect 14331 35404 14361 35438
rect 603 35396 14361 35404
rect 603 35370 807 35396
rect 603 35336 632 35370
rect 666 35362 807 35370
rect 841 35389 14361 35396
rect 841 35362 14122 35389
rect 666 35355 14122 35362
rect 14156 35370 14361 35389
rect 14156 35355 14297 35370
rect 666 35336 14297 35355
rect 14331 35336 14361 35370
rect 603 35324 14361 35336
rect 603 35302 807 35324
rect 603 35268 632 35302
rect 666 35290 807 35302
rect 841 35317 14361 35324
rect 841 35290 14122 35317
rect 666 35283 14122 35290
rect 14156 35302 14361 35317
rect 14156 35283 14297 35302
rect 666 35268 14297 35283
rect 14331 35268 14361 35302
rect 603 35252 14361 35268
rect 603 35234 807 35252
rect 603 35200 632 35234
rect 666 35218 807 35234
rect 841 35245 14361 35252
rect 841 35218 14122 35245
rect 666 35211 14122 35218
rect 14156 35234 14361 35245
rect 14156 35211 14297 35234
rect 666 35200 14297 35211
rect 14331 35200 14361 35234
rect 603 35180 14361 35200
rect 603 35166 807 35180
rect 603 35132 632 35166
rect 666 35146 807 35166
rect 841 35173 14361 35180
rect 841 35146 14122 35173
rect 666 35139 14122 35146
rect 14156 35166 14361 35173
rect 14156 35139 14297 35166
rect 666 35132 14297 35139
rect 14331 35132 14361 35166
rect 603 35108 14361 35132
rect 603 35098 807 35108
rect 603 35064 632 35098
rect 666 35074 807 35098
rect 841 35101 14361 35108
rect 841 35074 14122 35101
rect 666 35067 14122 35074
rect 14156 35098 14361 35101
rect 14156 35067 14297 35098
rect 666 35064 14297 35067
rect 14331 35064 14361 35098
rect 603 35036 14361 35064
rect 603 35030 807 35036
rect 603 34996 632 35030
rect 666 35002 807 35030
rect 841 35030 14361 35036
rect 841 35029 14297 35030
rect 841 35002 14122 35029
rect 666 34996 14122 35002
rect 603 34995 14122 34996
rect 14156 34996 14297 35029
rect 14331 34996 14361 35030
rect 14156 34995 14361 34996
rect 603 34964 14361 34995
rect 603 34962 807 34964
rect 603 34928 632 34962
rect 666 34930 807 34962
rect 841 34962 14361 34964
rect 841 34957 14297 34962
rect 841 34930 14122 34957
rect 666 34928 14122 34930
rect 603 34923 14122 34928
rect 14156 34928 14297 34957
rect 14331 34928 14361 34962
rect 14156 34923 14361 34928
rect 603 34894 14361 34923
rect 603 34860 632 34894
rect 666 34892 14297 34894
rect 666 34860 807 34892
rect 603 34858 807 34860
rect 841 34885 14297 34892
rect 841 34858 14122 34885
rect 603 34851 14122 34858
rect 14156 34860 14297 34885
rect 14331 34860 14361 34894
rect 14156 34851 14361 34860
rect 603 34831 14361 34851
rect 603 34826 1026 34831
rect 603 34792 632 34826
rect 666 34820 1026 34826
rect 666 34792 807 34820
rect 603 34786 807 34792
rect 841 34786 1026 34820
rect 603 34758 1026 34786
rect 603 34724 632 34758
rect 666 34748 1026 34758
rect 666 34724 807 34748
rect 603 34714 807 34724
rect 841 34714 1026 34748
rect 13968 34826 14361 34831
rect 13968 34813 14297 34826
rect 13968 34779 14122 34813
rect 14156 34792 14297 34813
rect 14331 34792 14361 34826
rect 14156 34779 14361 34792
rect 13968 34758 14361 34779
rect 13968 34741 14297 34758
rect 603 34690 1026 34714
rect 603 34656 632 34690
rect 666 34676 1026 34690
rect 666 34656 807 34676
rect 603 34642 807 34656
rect 841 34642 1026 34676
rect 603 34622 1026 34642
rect 603 34588 632 34622
rect 666 34604 1026 34622
rect 666 34588 807 34604
rect 603 34570 807 34588
rect 841 34570 1026 34604
rect 603 34554 1026 34570
rect 603 34520 632 34554
rect 666 34532 1026 34554
rect 666 34520 807 34532
rect 603 34498 807 34520
rect 841 34498 1026 34532
rect 603 34486 1026 34498
rect 603 34452 632 34486
rect 666 34460 1026 34486
rect 666 34452 807 34460
rect 603 34426 807 34452
rect 841 34426 1026 34460
rect 603 34418 1026 34426
rect 603 34384 632 34418
rect 666 34388 1026 34418
rect 666 34384 807 34388
rect 603 34354 807 34384
rect 841 34354 1026 34388
rect 603 34350 1026 34354
rect 603 34316 632 34350
rect 666 34316 1026 34350
rect 603 34282 807 34316
rect 841 34282 1026 34316
rect 603 34248 632 34282
rect 666 34248 1026 34282
rect 603 34244 1026 34248
rect 603 34214 807 34244
rect 603 34180 632 34214
rect 666 34210 807 34214
rect 841 34210 1026 34244
rect 666 34180 1026 34210
rect 603 34172 1026 34180
rect 603 34146 807 34172
rect 603 34112 632 34146
rect 666 34138 807 34146
rect 841 34138 1026 34172
rect 666 34112 1026 34138
rect 603 34100 1026 34112
rect 603 34078 807 34100
rect 603 34044 632 34078
rect 666 34066 807 34078
rect 841 34066 1026 34100
rect 666 34044 1026 34066
rect 603 34028 1026 34044
rect 603 34010 807 34028
rect 603 33976 632 34010
rect 666 33994 807 34010
rect 841 33994 1026 34028
rect 666 33976 1026 33994
rect 603 33956 1026 33976
rect 603 33942 807 33956
rect 603 33908 632 33942
rect 666 33922 807 33942
rect 841 33922 1026 33956
rect 666 33908 1026 33922
rect 603 33884 1026 33908
rect 603 33874 807 33884
rect 603 33840 632 33874
rect 666 33850 807 33874
rect 841 33850 1026 33884
rect 666 33840 1026 33850
rect 603 33812 1026 33840
rect 603 33806 807 33812
rect 603 33772 632 33806
rect 666 33778 807 33806
rect 841 33778 1026 33812
rect 666 33772 1026 33778
rect 603 33740 1026 33772
rect 603 33738 807 33740
rect 603 33704 632 33738
rect 666 33706 807 33738
rect 841 33706 1026 33740
rect 666 33704 1026 33706
rect 603 33670 1026 33704
rect 603 33636 632 33670
rect 666 33668 1026 33670
rect 666 33636 807 33668
rect 603 33634 807 33636
rect 841 33634 1026 33668
rect 603 33602 1026 33634
rect 603 33568 632 33602
rect 666 33596 1026 33602
rect 666 33568 807 33596
rect 603 33562 807 33568
rect 841 33562 1026 33596
rect 603 33534 1026 33562
rect 603 33500 632 33534
rect 666 33524 1026 33534
rect 666 33500 807 33524
rect 603 33490 807 33500
rect 841 33490 1026 33524
rect 603 33466 1026 33490
rect 603 33432 632 33466
rect 666 33452 1026 33466
rect 666 33432 807 33452
rect 603 33418 807 33432
rect 841 33418 1026 33452
rect 603 33398 1026 33418
rect 603 33364 632 33398
rect 666 33380 1026 33398
rect 666 33364 807 33380
rect 603 33346 807 33364
rect 841 33346 1026 33380
rect 603 33330 1026 33346
rect 603 33296 632 33330
rect 666 33308 1026 33330
rect 666 33296 807 33308
rect 603 33274 807 33296
rect 841 33274 1026 33308
rect 603 33262 1026 33274
rect 603 33228 632 33262
rect 666 33236 1026 33262
rect 666 33228 807 33236
rect 603 33202 807 33228
rect 841 33202 1026 33236
rect 603 33194 1026 33202
rect 603 33160 632 33194
rect 666 33164 1026 33194
rect 666 33160 807 33164
rect 603 33130 807 33160
rect 841 33130 1026 33164
rect 603 33126 1026 33130
rect 603 33092 632 33126
rect 666 33092 1026 33126
rect 603 33058 807 33092
rect 841 33058 1026 33092
rect 603 33024 632 33058
rect 666 33024 1026 33058
rect 603 33020 1026 33024
rect 603 32990 807 33020
rect 603 32956 632 32990
rect 666 32986 807 32990
rect 841 32986 1026 33020
rect 666 32956 1026 32986
rect 603 32948 1026 32956
rect 603 32922 807 32948
rect 603 32888 632 32922
rect 666 32914 807 32922
rect 841 32914 1026 32948
rect 666 32888 1026 32914
rect 603 32876 1026 32888
rect 603 32854 807 32876
rect 603 32820 632 32854
rect 666 32842 807 32854
rect 841 32842 1026 32876
rect 666 32820 1026 32842
rect 603 32804 1026 32820
rect 603 32786 807 32804
rect 603 32752 632 32786
rect 666 32770 807 32786
rect 841 32770 1026 32804
rect 666 32752 1026 32770
rect 603 32732 1026 32752
rect 603 32718 807 32732
rect 603 32684 632 32718
rect 666 32698 807 32718
rect 841 32698 1026 32732
rect 666 32684 1026 32698
rect 603 32660 1026 32684
rect 603 32650 807 32660
rect 603 32616 632 32650
rect 666 32626 807 32650
rect 841 32626 1026 32660
rect 666 32616 1026 32626
rect 603 32588 1026 32616
rect 603 32582 807 32588
rect 603 32548 632 32582
rect 666 32554 807 32582
rect 841 32554 1026 32588
rect 666 32548 1026 32554
rect 603 32516 1026 32548
rect 603 32514 807 32516
rect 603 32480 632 32514
rect 666 32482 807 32514
rect 841 32482 1026 32516
rect 666 32480 1026 32482
rect 603 32446 1026 32480
rect 603 32412 632 32446
rect 666 32444 1026 32446
rect 666 32412 807 32444
rect 603 32410 807 32412
rect 841 32410 1026 32444
rect 603 32378 1026 32410
rect 603 32344 632 32378
rect 666 32372 1026 32378
rect 666 32344 807 32372
rect 603 32338 807 32344
rect 841 32338 1026 32372
rect 603 32310 1026 32338
rect 603 32276 632 32310
rect 666 32300 1026 32310
rect 666 32276 807 32300
rect 603 32266 807 32276
rect 841 32266 1026 32300
rect 603 32242 1026 32266
rect 603 32208 632 32242
rect 666 32228 1026 32242
rect 666 32208 807 32228
rect 603 32194 807 32208
rect 841 32194 1026 32228
rect 603 32174 1026 32194
rect 603 32140 632 32174
rect 666 32156 1026 32174
rect 666 32140 807 32156
rect 603 32122 807 32140
rect 841 32122 1026 32156
rect 603 32106 1026 32122
rect 603 32072 632 32106
rect 666 32084 1026 32106
rect 666 32072 807 32084
rect 603 32050 807 32072
rect 841 32050 1026 32084
rect 603 32038 1026 32050
rect 603 32004 632 32038
rect 666 32012 1026 32038
rect 666 32004 807 32012
rect 603 31978 807 32004
rect 841 31978 1026 32012
rect 603 31970 1026 31978
rect 603 31936 632 31970
rect 666 31940 1026 31970
rect 666 31936 807 31940
rect 603 31906 807 31936
rect 841 31906 1026 31940
rect 603 31902 1026 31906
rect 603 31868 632 31902
rect 666 31868 1026 31902
rect 603 31834 807 31868
rect 841 31834 1026 31868
rect 603 31800 632 31834
rect 666 31800 1026 31834
rect 603 31796 1026 31800
rect 603 31766 807 31796
rect 603 31732 632 31766
rect 666 31762 807 31766
rect 841 31762 1026 31796
rect 666 31732 1026 31762
rect 603 31724 1026 31732
rect 603 31698 807 31724
rect 603 31664 632 31698
rect 666 31690 807 31698
rect 841 31690 1026 31724
rect 666 31664 1026 31690
rect 603 31652 1026 31664
rect 603 31630 807 31652
rect 603 31596 632 31630
rect 666 31618 807 31630
rect 841 31618 1026 31652
rect 666 31596 1026 31618
rect 603 31580 1026 31596
rect 603 31562 807 31580
rect 603 31528 632 31562
rect 666 31546 807 31562
rect 841 31546 1026 31580
rect 666 31528 1026 31546
rect 603 31508 1026 31528
rect 603 31494 807 31508
rect 603 31460 632 31494
rect 666 31474 807 31494
rect 841 31474 1026 31508
rect 666 31460 1026 31474
rect 603 31436 1026 31460
rect 603 31426 807 31436
rect 603 31392 632 31426
rect 666 31402 807 31426
rect 841 31402 1026 31436
rect 666 31392 1026 31402
rect 603 31364 1026 31392
rect 603 31358 807 31364
rect 603 31324 632 31358
rect 666 31330 807 31358
rect 841 31330 1026 31364
rect 666 31324 1026 31330
rect 603 31292 1026 31324
rect 603 31290 807 31292
rect 603 31256 632 31290
rect 666 31258 807 31290
rect 841 31258 1026 31292
rect 666 31256 1026 31258
rect 603 31222 1026 31256
rect 603 31188 632 31222
rect 666 31220 1026 31222
rect 666 31188 807 31220
rect 603 31186 807 31188
rect 841 31186 1026 31220
rect 603 31154 1026 31186
rect 603 31120 632 31154
rect 666 31148 1026 31154
rect 666 31120 807 31148
rect 603 31114 807 31120
rect 841 31114 1026 31148
rect 603 31086 1026 31114
rect 603 31052 632 31086
rect 666 31076 1026 31086
rect 666 31052 807 31076
rect 603 31042 807 31052
rect 841 31042 1026 31076
rect 603 31018 1026 31042
rect 603 30984 632 31018
rect 666 31004 1026 31018
rect 666 30984 807 31004
rect 603 30970 807 30984
rect 841 30970 1026 31004
rect 603 30950 1026 30970
rect 603 30916 632 30950
rect 666 30932 1026 30950
rect 666 30916 807 30932
rect 603 30898 807 30916
rect 841 30898 1026 30932
rect 603 30882 1026 30898
rect 603 30848 632 30882
rect 666 30860 1026 30882
rect 666 30848 807 30860
rect 603 30826 807 30848
rect 841 30826 1026 30860
rect 603 30814 1026 30826
rect 603 30780 632 30814
rect 666 30788 1026 30814
rect 666 30780 807 30788
rect 603 30754 807 30780
rect 841 30754 1026 30788
rect 603 30746 1026 30754
rect 603 30712 632 30746
rect 666 30716 1026 30746
rect 666 30712 807 30716
rect 603 30682 807 30712
rect 841 30682 1026 30716
rect 603 30678 1026 30682
rect 603 30644 632 30678
rect 666 30644 1026 30678
rect 603 30610 807 30644
rect 841 30610 1026 30644
rect 603 30576 632 30610
rect 666 30576 1026 30610
rect 603 30572 1026 30576
rect 603 30542 807 30572
rect 603 30508 632 30542
rect 666 30538 807 30542
rect 841 30538 1026 30572
rect 666 30508 1026 30538
rect 603 30500 1026 30508
rect 603 30474 807 30500
rect 603 30440 632 30474
rect 666 30466 807 30474
rect 841 30466 1026 30500
rect 666 30440 1026 30466
rect 603 30428 1026 30440
rect 603 30406 807 30428
rect 603 30372 632 30406
rect 666 30394 807 30406
rect 841 30394 1026 30428
rect 666 30372 1026 30394
rect 603 30356 1026 30372
rect 603 30338 807 30356
rect 603 30304 632 30338
rect 666 30322 807 30338
rect 841 30322 1026 30356
rect 666 30304 1026 30322
rect 603 30284 1026 30304
rect 603 30270 807 30284
rect 603 30236 632 30270
rect 666 30250 807 30270
rect 841 30250 1026 30284
rect 666 30236 1026 30250
rect 603 30212 1026 30236
rect 603 30202 807 30212
rect 603 30168 632 30202
rect 666 30178 807 30202
rect 841 30178 1026 30212
rect 666 30168 1026 30178
rect 603 30140 1026 30168
rect 603 30134 807 30140
rect 603 30100 632 30134
rect 666 30106 807 30134
rect 841 30106 1026 30140
rect 666 30100 1026 30106
rect 603 30068 1026 30100
rect 603 30066 807 30068
rect 603 30032 632 30066
rect 666 30034 807 30066
rect 841 30034 1026 30068
rect 666 30032 1026 30034
rect 603 29998 1026 30032
rect 603 29964 632 29998
rect 666 29996 1026 29998
rect 666 29964 807 29996
rect 603 29962 807 29964
rect 841 29962 1026 29996
rect 603 29930 1026 29962
rect 603 29896 632 29930
rect 666 29924 1026 29930
rect 666 29896 807 29924
rect 603 29890 807 29896
rect 841 29890 1026 29924
rect 603 29862 1026 29890
rect 603 29828 632 29862
rect 666 29852 1026 29862
rect 666 29828 807 29852
rect 603 29818 807 29828
rect 841 29818 1026 29852
rect 603 29794 1026 29818
rect 603 29760 632 29794
rect 666 29780 1026 29794
rect 666 29760 807 29780
rect 603 29746 807 29760
rect 841 29746 1026 29780
rect 603 29726 1026 29746
rect 603 29692 632 29726
rect 666 29708 1026 29726
rect 666 29692 807 29708
rect 603 29674 807 29692
rect 841 29674 1026 29708
rect 603 29658 1026 29674
rect 603 29624 632 29658
rect 666 29636 1026 29658
rect 666 29624 807 29636
rect 603 29602 807 29624
rect 841 29602 1026 29636
rect 603 29590 1026 29602
rect 603 29556 632 29590
rect 666 29564 1026 29590
rect 666 29556 807 29564
rect 603 29530 807 29556
rect 841 29530 1026 29564
rect 603 29522 1026 29530
rect 603 29488 632 29522
rect 666 29492 1026 29522
rect 666 29488 807 29492
rect 603 29458 807 29488
rect 841 29458 1026 29492
rect 603 29454 1026 29458
rect 603 29420 632 29454
rect 666 29420 1026 29454
rect 603 29386 807 29420
rect 841 29386 1026 29420
rect 603 29352 632 29386
rect 666 29352 1026 29386
rect 603 29348 1026 29352
rect 603 29318 807 29348
rect 603 29284 632 29318
rect 666 29314 807 29318
rect 841 29314 1026 29348
rect 666 29284 1026 29314
rect 603 29276 1026 29284
rect 603 29250 807 29276
rect 603 29216 632 29250
rect 666 29242 807 29250
rect 841 29242 1026 29276
rect 666 29216 1026 29242
rect 603 29204 1026 29216
rect 603 29182 807 29204
rect 603 29148 632 29182
rect 666 29170 807 29182
rect 841 29170 1026 29204
rect 666 29148 1026 29170
rect 603 29132 1026 29148
rect 603 29114 807 29132
rect 603 29080 632 29114
rect 666 29098 807 29114
rect 841 29098 1026 29132
rect 666 29080 1026 29098
rect 603 29060 1026 29080
rect 603 29046 807 29060
rect 603 29012 632 29046
rect 666 29026 807 29046
rect 841 29026 1026 29060
rect 666 29012 1026 29026
rect 603 28988 1026 29012
rect 603 28978 807 28988
rect 603 28944 632 28978
rect 666 28954 807 28978
rect 841 28954 1026 28988
rect 666 28944 1026 28954
rect 603 28916 1026 28944
rect 603 28910 807 28916
rect 603 28876 632 28910
rect 666 28882 807 28910
rect 841 28882 1026 28916
rect 666 28876 1026 28882
rect 603 28844 1026 28876
rect 603 28842 807 28844
rect 603 28808 632 28842
rect 666 28810 807 28842
rect 841 28810 1026 28844
rect 666 28808 1026 28810
rect 603 28774 1026 28808
rect 603 28740 632 28774
rect 666 28772 1026 28774
rect 666 28740 807 28772
rect 603 28738 807 28740
rect 841 28738 1026 28772
rect 603 28706 1026 28738
rect 603 28672 632 28706
rect 666 28700 1026 28706
rect 666 28672 807 28700
rect 603 28666 807 28672
rect 841 28666 1026 28700
rect 603 28638 1026 28666
rect 603 28604 632 28638
rect 666 28628 1026 28638
rect 666 28604 807 28628
rect 603 28594 807 28604
rect 841 28594 1026 28628
rect 603 28570 1026 28594
rect 603 28536 632 28570
rect 666 28556 1026 28570
rect 666 28536 807 28556
rect 603 28522 807 28536
rect 841 28522 1026 28556
rect 603 28502 1026 28522
rect 603 28468 632 28502
rect 666 28484 1026 28502
rect 666 28468 807 28484
rect 603 28450 807 28468
rect 841 28450 1026 28484
rect 603 28434 1026 28450
rect 603 28400 632 28434
rect 666 28412 1026 28434
rect 666 28400 807 28412
rect 603 28378 807 28400
rect 841 28378 1026 28412
rect 603 28366 1026 28378
rect 603 28332 632 28366
rect 666 28340 1026 28366
rect 666 28332 807 28340
rect 603 28306 807 28332
rect 841 28306 1026 28340
rect 603 28298 1026 28306
rect 603 28264 632 28298
rect 666 28268 1026 28298
rect 666 28264 807 28268
rect 603 28234 807 28264
rect 841 28234 1026 28268
rect 603 28230 1026 28234
rect 603 28196 632 28230
rect 666 28196 1026 28230
rect 603 28162 807 28196
rect 841 28162 1026 28196
rect 603 28128 632 28162
rect 666 28128 1026 28162
rect 603 28124 1026 28128
rect 603 28094 807 28124
rect 603 28060 632 28094
rect 666 28090 807 28094
rect 841 28090 1026 28124
rect 666 28060 1026 28090
rect 603 28052 1026 28060
rect 603 28026 807 28052
rect 603 27992 632 28026
rect 666 28018 807 28026
rect 841 28018 1026 28052
rect 666 27992 1026 28018
rect 603 27980 1026 27992
rect 603 27958 807 27980
rect 603 27924 632 27958
rect 666 27946 807 27958
rect 841 27946 1026 27980
rect 666 27924 1026 27946
rect 603 27908 1026 27924
rect 603 27890 807 27908
rect 603 27856 632 27890
rect 666 27874 807 27890
rect 841 27874 1026 27908
rect 666 27856 1026 27874
rect 603 27836 1026 27856
rect 603 27822 807 27836
rect 603 27788 632 27822
rect 666 27802 807 27822
rect 841 27802 1026 27836
rect 666 27788 1026 27802
rect 603 27764 1026 27788
rect 603 27754 807 27764
rect 603 27720 632 27754
rect 666 27730 807 27754
rect 841 27730 1026 27764
rect 666 27720 1026 27730
rect 603 27692 1026 27720
rect 603 27686 807 27692
rect 603 27652 632 27686
rect 666 27658 807 27686
rect 841 27658 1026 27692
rect 666 27652 1026 27658
rect 603 27620 1026 27652
rect 603 27618 807 27620
rect 603 27584 632 27618
rect 666 27586 807 27618
rect 841 27586 1026 27620
rect 666 27584 1026 27586
rect 603 27550 1026 27584
rect 603 27516 632 27550
rect 666 27548 1026 27550
rect 666 27516 807 27548
rect 603 27514 807 27516
rect 841 27514 1026 27548
rect 603 27482 1026 27514
rect 603 27448 632 27482
rect 666 27476 1026 27482
rect 666 27448 807 27476
rect 603 27442 807 27448
rect 841 27442 1026 27476
rect 603 27414 1026 27442
rect 603 27380 632 27414
rect 666 27404 1026 27414
rect 666 27380 807 27404
rect 603 27370 807 27380
rect 841 27370 1026 27404
rect 603 27346 1026 27370
rect 603 27312 632 27346
rect 666 27332 1026 27346
rect 666 27312 807 27332
rect 603 27298 807 27312
rect 841 27298 1026 27332
rect 603 27278 1026 27298
rect 603 27244 632 27278
rect 666 27260 1026 27278
rect 666 27244 807 27260
rect 603 27226 807 27244
rect 841 27226 1026 27260
rect 603 27210 1026 27226
rect 603 27176 632 27210
rect 666 27188 1026 27210
rect 666 27176 807 27188
rect 603 27154 807 27176
rect 841 27154 1026 27188
rect 603 27142 1026 27154
rect 603 27108 632 27142
rect 666 27116 1026 27142
rect 666 27108 807 27116
rect 603 27082 807 27108
rect 841 27082 1026 27116
rect 603 27074 1026 27082
rect 603 27040 632 27074
rect 666 27044 1026 27074
rect 666 27040 807 27044
rect 603 27010 807 27040
rect 841 27010 1026 27044
rect 603 27006 1026 27010
rect 603 26972 632 27006
rect 666 26972 1026 27006
rect 603 26938 807 26972
rect 841 26938 1026 26972
rect 603 26904 632 26938
rect 666 26904 1026 26938
rect 603 26900 1026 26904
rect 603 26870 807 26900
rect 603 26836 632 26870
rect 666 26866 807 26870
rect 841 26866 1026 26900
rect 666 26836 1026 26866
rect 603 26828 1026 26836
rect 603 26802 807 26828
rect 603 26768 632 26802
rect 666 26794 807 26802
rect 841 26794 1026 26828
rect 666 26768 1026 26794
rect 603 26756 1026 26768
rect 603 26734 807 26756
rect 603 26700 632 26734
rect 666 26722 807 26734
rect 841 26722 1026 26756
rect 666 26700 1026 26722
rect 603 26684 1026 26700
rect 603 26666 807 26684
rect 603 26632 632 26666
rect 666 26650 807 26666
rect 841 26650 1026 26684
rect 666 26632 1026 26650
rect 603 26612 1026 26632
rect 603 26598 807 26612
rect 603 26564 632 26598
rect 666 26578 807 26598
rect 841 26578 1026 26612
rect 666 26564 1026 26578
rect 603 26540 1026 26564
rect 603 26530 807 26540
rect 603 26496 632 26530
rect 666 26506 807 26530
rect 841 26506 1026 26540
rect 666 26496 1026 26506
rect 603 26468 1026 26496
rect 603 26462 807 26468
rect 603 26428 632 26462
rect 666 26434 807 26462
rect 841 26434 1026 26468
rect 666 26428 1026 26434
rect 603 26396 1026 26428
rect 603 26394 807 26396
rect 603 26360 632 26394
rect 666 26362 807 26394
rect 841 26362 1026 26396
rect 666 26360 1026 26362
rect 603 26326 1026 26360
rect 603 26292 632 26326
rect 666 26324 1026 26326
rect 666 26292 807 26324
rect 603 26290 807 26292
rect 841 26290 1026 26324
rect 603 26258 1026 26290
rect 603 26224 632 26258
rect 666 26252 1026 26258
rect 666 26224 807 26252
rect 603 26218 807 26224
rect 841 26218 1026 26252
rect 603 26190 1026 26218
rect 603 26156 632 26190
rect 666 26180 1026 26190
rect 666 26156 807 26180
rect 603 26146 807 26156
rect 841 26146 1026 26180
rect 603 26122 1026 26146
rect 603 26088 632 26122
rect 666 26108 1026 26122
rect 666 26088 807 26108
rect 603 26074 807 26088
rect 841 26074 1026 26108
rect 603 26054 1026 26074
rect 603 26020 632 26054
rect 666 26036 1026 26054
rect 666 26020 807 26036
rect 603 26002 807 26020
rect 841 26002 1026 26036
rect 603 25986 1026 26002
rect 603 25952 632 25986
rect 666 25964 1026 25986
rect 666 25952 807 25964
rect 603 25930 807 25952
rect 841 25930 1026 25964
rect 603 25918 1026 25930
rect 603 25884 632 25918
rect 666 25892 1026 25918
rect 666 25884 807 25892
rect 603 25858 807 25884
rect 841 25858 1026 25892
rect 603 25850 1026 25858
rect 603 25816 632 25850
rect 666 25820 1026 25850
rect 666 25816 807 25820
rect 603 25786 807 25816
rect 841 25786 1026 25820
rect 603 25782 1026 25786
rect 603 25748 632 25782
rect 666 25748 1026 25782
rect 603 25714 807 25748
rect 841 25714 1026 25748
rect 603 25680 632 25714
rect 666 25680 1026 25714
rect 603 25676 1026 25680
rect 603 25646 807 25676
rect 603 25612 632 25646
rect 666 25642 807 25646
rect 841 25642 1026 25676
rect 666 25612 1026 25642
rect 603 25604 1026 25612
rect 603 25578 807 25604
rect 603 25544 632 25578
rect 666 25570 807 25578
rect 841 25570 1026 25604
rect 666 25544 1026 25570
rect 603 25532 1026 25544
rect 603 25510 807 25532
rect 603 25476 632 25510
rect 666 25498 807 25510
rect 841 25498 1026 25532
rect 666 25476 1026 25498
rect 603 25460 1026 25476
rect 603 25442 807 25460
rect 603 25408 632 25442
rect 666 25426 807 25442
rect 841 25426 1026 25460
rect 666 25408 1026 25426
rect 603 25388 1026 25408
rect 603 25374 807 25388
rect 603 25340 632 25374
rect 666 25354 807 25374
rect 841 25354 1026 25388
rect 666 25340 1026 25354
rect 603 25316 1026 25340
rect 603 25306 807 25316
rect 603 25272 632 25306
rect 666 25282 807 25306
rect 841 25282 1026 25316
rect 666 25272 1026 25282
rect 603 25244 1026 25272
rect 603 25238 807 25244
rect 603 25204 632 25238
rect 666 25210 807 25238
rect 841 25210 1026 25244
rect 666 25204 1026 25210
rect 603 25172 1026 25204
rect 603 25170 807 25172
rect 603 25136 632 25170
rect 666 25138 807 25170
rect 841 25138 1026 25172
rect 666 25136 1026 25138
rect 603 25102 1026 25136
rect 603 25068 632 25102
rect 666 25100 1026 25102
rect 666 25068 807 25100
rect 603 25066 807 25068
rect 841 25066 1026 25100
rect 603 25034 1026 25066
rect 603 25000 632 25034
rect 666 25028 1026 25034
rect 666 25000 807 25028
rect 603 24994 807 25000
rect 841 24994 1026 25028
rect 603 24966 1026 24994
rect 603 24932 632 24966
rect 666 24956 1026 24966
rect 666 24932 807 24956
rect 603 24922 807 24932
rect 841 24922 1026 24956
rect 603 24898 1026 24922
rect 603 24864 632 24898
rect 666 24884 1026 24898
rect 666 24864 807 24884
rect 603 24850 807 24864
rect 841 24850 1026 24884
rect 603 24830 1026 24850
rect 603 24796 632 24830
rect 666 24812 1026 24830
rect 666 24796 807 24812
rect 603 24778 807 24796
rect 841 24778 1026 24812
rect 603 24762 1026 24778
rect 603 24728 632 24762
rect 666 24740 1026 24762
rect 666 24728 807 24740
rect 603 24706 807 24728
rect 841 24706 1026 24740
rect 603 24694 1026 24706
rect 603 24660 632 24694
rect 666 24668 1026 24694
rect 666 24660 807 24668
rect 603 24634 807 24660
rect 841 24634 1026 24668
rect 603 24626 1026 24634
rect 603 24592 632 24626
rect 666 24596 1026 24626
rect 666 24592 807 24596
rect 603 24562 807 24592
rect 841 24562 1026 24596
rect 603 24558 1026 24562
rect 603 24524 632 24558
rect 666 24524 1026 24558
rect 603 24490 807 24524
rect 841 24490 1026 24524
rect 603 24456 632 24490
rect 666 24456 1026 24490
rect 603 24452 1026 24456
rect 603 24422 807 24452
rect 603 24388 632 24422
rect 666 24418 807 24422
rect 841 24418 1026 24452
rect 666 24388 1026 24418
rect 603 24380 1026 24388
rect 603 24354 807 24380
rect 603 24320 632 24354
rect 666 24346 807 24354
rect 841 24346 1026 24380
rect 666 24320 1026 24346
rect 603 24308 1026 24320
rect 603 24286 807 24308
rect 603 24252 632 24286
rect 666 24274 807 24286
rect 841 24274 1026 24308
rect 666 24252 1026 24274
rect 603 24236 1026 24252
rect 603 24218 807 24236
rect 603 24184 632 24218
rect 666 24202 807 24218
rect 841 24202 1026 24236
rect 666 24184 1026 24202
rect 603 24164 1026 24184
rect 603 24150 807 24164
rect 603 24116 632 24150
rect 666 24130 807 24150
rect 841 24130 1026 24164
rect 666 24116 1026 24130
rect 603 24092 1026 24116
rect 603 24082 807 24092
rect 603 24048 632 24082
rect 666 24058 807 24082
rect 841 24058 1026 24092
rect 666 24048 1026 24058
rect 603 24020 1026 24048
rect 603 24014 807 24020
rect 603 23980 632 24014
rect 666 23986 807 24014
rect 841 23986 1026 24020
rect 666 23980 1026 23986
rect 603 23948 1026 23980
rect 603 23946 807 23948
rect 603 23912 632 23946
rect 666 23914 807 23946
rect 841 23914 1026 23948
rect 666 23912 1026 23914
rect 603 23878 1026 23912
rect 603 23844 632 23878
rect 666 23876 1026 23878
rect 666 23844 807 23876
rect 603 23842 807 23844
rect 841 23842 1026 23876
rect 603 23810 1026 23842
rect 603 23776 632 23810
rect 666 23804 1026 23810
rect 666 23776 807 23804
rect 603 23770 807 23776
rect 841 23770 1026 23804
rect 603 23742 1026 23770
rect 603 23708 632 23742
rect 666 23732 1026 23742
rect 666 23708 807 23732
rect 603 23698 807 23708
rect 841 23698 1026 23732
rect 603 23674 1026 23698
rect 603 23640 632 23674
rect 666 23660 1026 23674
rect 666 23640 807 23660
rect 603 23626 807 23640
rect 841 23626 1026 23660
rect 603 23606 1026 23626
rect 603 23572 632 23606
rect 666 23588 1026 23606
rect 666 23572 807 23588
rect 603 23554 807 23572
rect 841 23554 1026 23588
rect 603 23538 1026 23554
rect 603 23504 632 23538
rect 666 23516 1026 23538
rect 666 23504 807 23516
rect 603 23482 807 23504
rect 841 23482 1026 23516
rect 603 23470 1026 23482
rect 603 23436 632 23470
rect 666 23444 1026 23470
rect 666 23436 807 23444
rect 603 23410 807 23436
rect 841 23410 1026 23444
rect 603 23402 1026 23410
rect 603 23368 632 23402
rect 666 23372 1026 23402
rect 666 23368 807 23372
rect 603 23338 807 23368
rect 841 23338 1026 23372
rect 603 23334 1026 23338
rect 603 23300 632 23334
rect 666 23300 1026 23334
rect 603 23266 807 23300
rect 841 23266 1026 23300
rect 603 23232 632 23266
rect 666 23232 1026 23266
rect 603 23228 1026 23232
rect 603 23198 807 23228
rect 603 23164 632 23198
rect 666 23194 807 23198
rect 841 23194 1026 23228
rect 666 23164 1026 23194
rect 603 23156 1026 23164
rect 603 23130 807 23156
rect 603 23096 632 23130
rect 666 23122 807 23130
rect 841 23122 1026 23156
rect 666 23096 1026 23122
rect 603 23084 1026 23096
rect 603 23062 807 23084
rect 603 23028 632 23062
rect 666 23050 807 23062
rect 841 23050 1026 23084
rect 666 23028 1026 23050
rect 603 23012 1026 23028
rect 603 22994 807 23012
rect 603 22960 632 22994
rect 666 22978 807 22994
rect 841 22978 1026 23012
rect 666 22960 1026 22978
rect 603 22940 1026 22960
rect 603 22926 807 22940
rect 603 22892 632 22926
rect 666 22906 807 22926
rect 841 22906 1026 22940
rect 666 22892 1026 22906
rect 603 22868 1026 22892
rect 603 22858 807 22868
rect 603 22824 632 22858
rect 666 22834 807 22858
rect 841 22834 1026 22868
rect 666 22824 1026 22834
rect 603 22796 1026 22824
rect 603 22790 807 22796
rect 603 22756 632 22790
rect 666 22762 807 22790
rect 841 22762 1026 22796
rect 666 22756 1026 22762
rect 603 22724 1026 22756
rect 603 22722 807 22724
rect 603 22688 632 22722
rect 666 22690 807 22722
rect 841 22690 1026 22724
rect 666 22688 1026 22690
rect 603 22654 1026 22688
rect 603 22620 632 22654
rect 666 22652 1026 22654
rect 666 22620 807 22652
rect 603 22618 807 22620
rect 841 22618 1026 22652
rect 603 22586 1026 22618
rect 603 22552 632 22586
rect 666 22580 1026 22586
rect 666 22552 807 22580
rect 603 22546 807 22552
rect 841 22546 1026 22580
rect 603 22518 1026 22546
rect 603 22484 632 22518
rect 666 22508 1026 22518
rect 666 22484 807 22508
rect 603 22474 807 22484
rect 841 22474 1026 22508
rect 603 22450 1026 22474
rect 603 22416 632 22450
rect 666 22436 1026 22450
rect 666 22416 807 22436
rect 603 22402 807 22416
rect 841 22402 1026 22436
rect 603 22382 1026 22402
rect 603 22348 632 22382
rect 666 22364 1026 22382
rect 666 22348 807 22364
rect 603 22330 807 22348
rect 841 22330 1026 22364
rect 603 22314 1026 22330
rect 603 22280 632 22314
rect 666 22292 1026 22314
rect 666 22280 807 22292
rect 603 22258 807 22280
rect 841 22258 1026 22292
rect 603 22246 1026 22258
rect 603 22212 632 22246
rect 666 22220 1026 22246
rect 666 22212 807 22220
rect 603 22186 807 22212
rect 841 22186 1026 22220
rect 603 22178 1026 22186
rect 603 22144 632 22178
rect 666 22148 1026 22178
rect 666 22144 807 22148
rect 603 22114 807 22144
rect 841 22114 1026 22148
rect 603 22110 1026 22114
rect 603 22076 632 22110
rect 666 22076 1026 22110
rect 603 22042 807 22076
rect 841 22042 1026 22076
rect 603 22008 632 22042
rect 666 22008 1026 22042
rect 603 22004 1026 22008
rect 603 21974 807 22004
rect 603 21940 632 21974
rect 666 21970 807 21974
rect 841 21970 1026 22004
rect 666 21940 1026 21970
rect 603 21932 1026 21940
rect 603 21906 807 21932
rect 603 21872 632 21906
rect 666 21898 807 21906
rect 841 21898 1026 21932
rect 666 21872 1026 21898
rect 603 21860 1026 21872
rect 603 21838 807 21860
rect 603 21804 632 21838
rect 666 21826 807 21838
rect 841 21826 1026 21860
rect 666 21804 1026 21826
rect 603 21788 1026 21804
rect 603 21770 807 21788
rect 603 21736 632 21770
rect 666 21754 807 21770
rect 841 21754 1026 21788
rect 666 21736 1026 21754
rect 603 21716 1026 21736
rect 603 21702 807 21716
rect 603 21668 632 21702
rect 666 21682 807 21702
rect 841 21682 1026 21716
rect 666 21668 1026 21682
rect 603 21644 1026 21668
rect 603 21634 807 21644
rect 603 21600 632 21634
rect 666 21610 807 21634
rect 841 21610 1026 21644
rect 666 21600 1026 21610
rect 603 21572 1026 21600
rect 603 21566 807 21572
rect 603 21532 632 21566
rect 666 21538 807 21566
rect 841 21538 1026 21572
rect 666 21532 1026 21538
rect 603 21500 1026 21532
rect 603 21498 807 21500
rect 603 21464 632 21498
rect 666 21466 807 21498
rect 841 21466 1026 21500
rect 666 21464 1026 21466
rect 603 21430 1026 21464
rect 603 21396 632 21430
rect 666 21428 1026 21430
rect 666 21396 807 21428
rect 603 21394 807 21396
rect 841 21394 1026 21428
rect 603 21362 1026 21394
rect 603 21328 632 21362
rect 666 21356 1026 21362
rect 666 21328 807 21356
rect 603 21322 807 21328
rect 841 21322 1026 21356
rect 603 21294 1026 21322
rect 603 21260 632 21294
rect 666 21284 1026 21294
rect 666 21260 807 21284
rect 603 21250 807 21260
rect 841 21250 1026 21284
rect 603 21226 1026 21250
rect 603 21192 632 21226
rect 666 21212 1026 21226
rect 666 21192 807 21212
rect 603 21178 807 21192
rect 841 21178 1026 21212
rect 603 21158 1026 21178
rect 603 21124 632 21158
rect 666 21140 1026 21158
rect 666 21124 807 21140
rect 603 21106 807 21124
rect 841 21106 1026 21140
rect 603 21090 1026 21106
rect 603 21056 632 21090
rect 666 21068 1026 21090
rect 666 21056 807 21068
rect 603 21034 807 21056
rect 841 21034 1026 21068
rect 603 21022 1026 21034
rect 603 20988 632 21022
rect 666 20996 1026 21022
rect 666 20988 807 20996
rect 603 20962 807 20988
rect 841 20962 1026 20996
rect 603 20954 1026 20962
rect 603 20920 632 20954
rect 666 20924 1026 20954
rect 666 20920 807 20924
rect 603 20890 807 20920
rect 841 20890 1026 20924
rect 603 20886 1026 20890
rect 603 20852 632 20886
rect 666 20852 1026 20886
rect 603 20818 807 20852
rect 841 20818 1026 20852
rect 603 20784 632 20818
rect 666 20784 1026 20818
rect 603 20780 1026 20784
rect 603 20750 807 20780
rect 603 20716 632 20750
rect 666 20746 807 20750
rect 841 20746 1026 20780
rect 666 20716 1026 20746
rect 603 20708 1026 20716
rect 603 20682 807 20708
rect 603 20648 632 20682
rect 666 20674 807 20682
rect 841 20674 1026 20708
rect 666 20648 1026 20674
rect 603 20636 1026 20648
rect 603 20614 807 20636
rect 603 20580 632 20614
rect 666 20602 807 20614
rect 841 20602 1026 20636
rect 666 20580 1026 20602
rect 603 20564 1026 20580
rect 603 20546 807 20564
rect 603 20512 632 20546
rect 666 20530 807 20546
rect 841 20530 1026 20564
rect 666 20512 1026 20530
rect 603 20492 1026 20512
rect 603 20478 807 20492
rect 603 20444 632 20478
rect 666 20458 807 20478
rect 841 20458 1026 20492
rect 666 20444 1026 20458
rect 603 20420 1026 20444
rect 603 20410 807 20420
rect 603 20376 632 20410
rect 666 20386 807 20410
rect 841 20386 1026 20420
rect 666 20376 1026 20386
rect 603 20348 1026 20376
rect 603 20342 807 20348
rect 603 20308 632 20342
rect 666 20314 807 20342
rect 841 20314 1026 20348
rect 666 20308 1026 20314
rect 603 20276 1026 20308
rect 603 20274 807 20276
rect 603 20240 632 20274
rect 666 20242 807 20274
rect 841 20242 1026 20276
rect 666 20240 1026 20242
rect 603 20206 1026 20240
rect 603 20172 632 20206
rect 666 20204 1026 20206
rect 666 20172 807 20204
rect 603 20170 807 20172
rect 841 20170 1026 20204
rect 603 20138 1026 20170
rect 603 20104 632 20138
rect 666 20132 1026 20138
rect 666 20104 807 20132
rect 603 20098 807 20104
rect 841 20098 1026 20132
rect 603 20070 1026 20098
rect 603 20036 632 20070
rect 666 20060 1026 20070
rect 666 20036 807 20060
rect 603 20026 807 20036
rect 841 20026 1026 20060
rect 603 20002 1026 20026
rect 603 19968 632 20002
rect 666 19988 1026 20002
rect 666 19968 807 19988
rect 603 19954 807 19968
rect 841 19954 1026 19988
rect 603 19934 1026 19954
rect 603 19900 632 19934
rect 666 19916 1026 19934
rect 666 19900 807 19916
rect 603 19882 807 19900
rect 841 19882 1026 19916
rect 603 19866 1026 19882
rect 603 19832 632 19866
rect 666 19844 1026 19866
rect 666 19832 807 19844
rect 603 19810 807 19832
rect 841 19810 1026 19844
rect 603 19798 1026 19810
rect 603 19764 632 19798
rect 666 19772 1026 19798
rect 666 19764 807 19772
rect 603 19738 807 19764
rect 841 19738 1026 19772
rect 603 19730 1026 19738
rect 603 19696 632 19730
rect 666 19700 1026 19730
rect 666 19696 807 19700
rect 603 19666 807 19696
rect 841 19666 1026 19700
rect 603 19662 1026 19666
rect 603 19628 632 19662
rect 666 19628 1026 19662
rect 603 19594 807 19628
rect 841 19594 1026 19628
rect 603 19560 632 19594
rect 666 19560 1026 19594
rect 603 19556 1026 19560
rect 603 19526 807 19556
rect 603 19492 632 19526
rect 666 19522 807 19526
rect 841 19522 1026 19556
rect 666 19492 1026 19522
rect 603 19484 1026 19492
rect 603 19458 807 19484
rect 603 19424 632 19458
rect 666 19450 807 19458
rect 841 19450 1026 19484
rect 666 19424 1026 19450
rect 603 19412 1026 19424
rect 603 19390 807 19412
rect 603 19356 632 19390
rect 666 19378 807 19390
rect 841 19378 1026 19412
rect 666 19356 1026 19378
rect 603 19340 1026 19356
rect 603 19322 807 19340
rect 603 19288 632 19322
rect 666 19306 807 19322
rect 841 19306 1026 19340
rect 666 19288 1026 19306
rect 603 19268 1026 19288
rect 603 19254 807 19268
rect 603 19220 632 19254
rect 666 19234 807 19254
rect 841 19234 1026 19268
rect 666 19220 1026 19234
rect 603 19196 1026 19220
rect 603 19186 807 19196
rect 603 19152 632 19186
rect 666 19162 807 19186
rect 841 19162 1026 19196
rect 666 19152 1026 19162
rect 603 19124 1026 19152
rect 603 19118 807 19124
rect 603 19084 632 19118
rect 666 19090 807 19118
rect 841 19090 1026 19124
rect 666 19084 1026 19090
rect 603 19052 1026 19084
rect 603 19050 807 19052
rect 603 19016 632 19050
rect 666 19018 807 19050
rect 841 19018 1026 19052
rect 666 19016 1026 19018
rect 603 18982 1026 19016
rect 603 18948 632 18982
rect 666 18980 1026 18982
rect 666 18948 807 18980
rect 603 18946 807 18948
rect 841 18946 1026 18980
rect 603 18914 1026 18946
rect 603 18880 632 18914
rect 666 18908 1026 18914
rect 666 18880 807 18908
rect 603 18874 807 18880
rect 841 18874 1026 18908
rect 603 18846 1026 18874
rect 603 18812 632 18846
rect 666 18836 1026 18846
rect 666 18812 807 18836
rect 603 18802 807 18812
rect 841 18802 1026 18836
rect 603 18778 1026 18802
rect 603 18744 632 18778
rect 666 18764 1026 18778
rect 666 18744 807 18764
rect 603 18730 807 18744
rect 841 18730 1026 18764
rect 603 18710 1026 18730
rect 603 18676 632 18710
rect 666 18692 1026 18710
rect 666 18676 807 18692
rect 603 18658 807 18676
rect 841 18658 1026 18692
rect 603 18642 1026 18658
rect 603 18608 632 18642
rect 666 18620 1026 18642
rect 666 18608 807 18620
rect 603 18586 807 18608
rect 841 18586 1026 18620
rect 603 18574 1026 18586
rect 603 18540 632 18574
rect 666 18548 1026 18574
rect 666 18540 807 18548
rect 603 18514 807 18540
rect 841 18514 1026 18548
rect 603 18506 1026 18514
rect 603 18472 632 18506
rect 666 18476 1026 18506
rect 666 18472 807 18476
rect 603 18442 807 18472
rect 841 18442 1026 18476
rect 603 18438 1026 18442
rect 603 18404 632 18438
rect 666 18404 1026 18438
rect 603 18370 807 18404
rect 841 18370 1026 18404
rect 603 18336 632 18370
rect 666 18336 1026 18370
rect 603 18332 1026 18336
rect 603 18302 807 18332
rect 603 18268 632 18302
rect 666 18298 807 18302
rect 841 18298 1026 18332
rect 666 18268 1026 18298
rect 603 18260 1026 18268
rect 603 18234 807 18260
rect 603 18200 632 18234
rect 666 18226 807 18234
rect 841 18226 1026 18260
rect 666 18200 1026 18226
rect 603 18188 1026 18200
rect 603 18166 807 18188
rect 603 18132 632 18166
rect 666 18154 807 18166
rect 841 18154 1026 18188
rect 666 18132 1026 18154
rect 603 18116 1026 18132
rect 603 18098 807 18116
rect 603 18064 632 18098
rect 666 18082 807 18098
rect 841 18082 1026 18116
rect 666 18064 1026 18082
rect 603 18044 1026 18064
rect 603 18030 807 18044
rect 603 17996 632 18030
rect 666 18010 807 18030
rect 841 18010 1026 18044
rect 666 17996 1026 18010
rect 603 17972 1026 17996
rect 603 17962 807 17972
rect 603 17928 632 17962
rect 666 17938 807 17962
rect 841 17938 1026 17972
rect 666 17928 1026 17938
rect 603 17900 1026 17928
rect 603 17894 807 17900
rect 603 17860 632 17894
rect 666 17866 807 17894
rect 841 17866 1026 17900
rect 666 17860 1026 17866
rect 603 17828 1026 17860
rect 603 17826 807 17828
rect 603 17792 632 17826
rect 666 17794 807 17826
rect 841 17794 1026 17828
rect 666 17792 1026 17794
rect 603 17758 1026 17792
rect 603 17724 632 17758
rect 666 17756 1026 17758
rect 666 17724 807 17756
rect 603 17722 807 17724
rect 841 17722 1026 17756
rect 603 17690 1026 17722
rect 603 17656 632 17690
rect 666 17684 1026 17690
rect 666 17656 807 17684
rect 603 17650 807 17656
rect 841 17650 1026 17684
rect 603 17622 1026 17650
rect 603 17588 632 17622
rect 666 17612 1026 17622
rect 666 17588 807 17612
rect 603 17578 807 17588
rect 841 17578 1026 17612
rect 603 17554 1026 17578
rect 603 17520 632 17554
rect 666 17540 1026 17554
rect 666 17520 807 17540
rect 603 17506 807 17520
rect 841 17506 1026 17540
rect 603 17486 1026 17506
rect 603 17452 632 17486
rect 666 17468 1026 17486
rect 666 17452 807 17468
rect 603 17434 807 17452
rect 841 17434 1026 17468
rect 603 17418 1026 17434
rect 603 17384 632 17418
rect 666 17396 1026 17418
rect 666 17384 807 17396
rect 603 17362 807 17384
rect 841 17362 1026 17396
rect 603 17350 1026 17362
rect 603 17316 632 17350
rect 666 17324 1026 17350
rect 666 17316 807 17324
rect 603 17290 807 17316
rect 841 17290 1026 17324
rect 603 17282 1026 17290
rect 603 17248 632 17282
rect 666 17252 1026 17282
rect 666 17248 807 17252
rect 603 17218 807 17248
rect 841 17218 1026 17252
rect 603 17214 1026 17218
rect 603 17180 632 17214
rect 666 17180 1026 17214
rect 603 17146 807 17180
rect 841 17146 1026 17180
rect 603 17112 632 17146
rect 666 17112 1026 17146
rect 603 17108 1026 17112
rect 603 17078 807 17108
rect 603 17044 632 17078
rect 666 17074 807 17078
rect 841 17074 1026 17108
rect 666 17044 1026 17074
rect 603 17036 1026 17044
rect 603 17010 807 17036
rect 603 16976 632 17010
rect 666 17002 807 17010
rect 841 17002 1026 17036
rect 666 16976 1026 17002
rect 603 16964 1026 16976
rect 603 16942 807 16964
rect 603 16908 632 16942
rect 666 16930 807 16942
rect 841 16930 1026 16964
rect 666 16908 1026 16930
rect 603 16892 1026 16908
rect 603 16874 807 16892
rect 603 16840 632 16874
rect 666 16858 807 16874
rect 841 16858 1026 16892
rect 666 16840 1026 16858
rect 603 16820 1026 16840
rect 603 16806 807 16820
rect 603 16772 632 16806
rect 666 16786 807 16806
rect 841 16786 1026 16820
rect 666 16772 1026 16786
rect 603 16748 1026 16772
rect 603 16738 807 16748
rect 603 16704 632 16738
rect 666 16714 807 16738
rect 841 16714 1026 16748
rect 666 16704 1026 16714
rect 603 16676 1026 16704
rect 603 16670 807 16676
rect 603 16636 632 16670
rect 666 16642 807 16670
rect 841 16642 1026 16676
rect 666 16636 1026 16642
rect 603 16604 1026 16636
rect 603 16602 807 16604
rect 603 16568 632 16602
rect 666 16570 807 16602
rect 841 16570 1026 16604
rect 666 16568 1026 16570
rect 603 16534 1026 16568
rect 603 16500 632 16534
rect 666 16532 1026 16534
rect 666 16500 807 16532
rect 603 16498 807 16500
rect 841 16498 1026 16532
rect 603 16466 1026 16498
rect 603 16432 632 16466
rect 666 16460 1026 16466
rect 666 16432 807 16460
rect 603 16426 807 16432
rect 841 16426 1026 16460
rect 603 16398 1026 16426
rect 603 16364 632 16398
rect 666 16388 1026 16398
rect 666 16364 807 16388
rect 603 16354 807 16364
rect 841 16354 1026 16388
rect 603 16330 1026 16354
rect 603 16296 632 16330
rect 666 16316 1026 16330
rect 666 16296 807 16316
rect 603 16282 807 16296
rect 841 16282 1026 16316
rect 603 16262 1026 16282
rect 603 16228 632 16262
rect 666 16244 1026 16262
rect 666 16228 807 16244
rect 603 16210 807 16228
rect 841 16210 1026 16244
rect 603 16194 1026 16210
rect 603 16160 632 16194
rect 666 16172 1026 16194
rect 666 16160 807 16172
rect 603 16138 807 16160
rect 841 16138 1026 16172
rect 603 16126 1026 16138
rect 603 16092 632 16126
rect 666 16100 1026 16126
rect 666 16092 807 16100
rect 603 16066 807 16092
rect 841 16066 1026 16100
rect 603 16058 1026 16066
rect 603 16024 632 16058
rect 666 16028 1026 16058
rect 666 16024 807 16028
rect 603 15994 807 16024
rect 841 15994 1026 16028
rect 603 15990 1026 15994
rect 603 15956 632 15990
rect 666 15956 1026 15990
rect 603 15922 807 15956
rect 841 15922 1026 15956
rect 603 15888 632 15922
rect 666 15888 1026 15922
rect 603 15884 1026 15888
rect 603 15854 807 15884
rect 603 15820 632 15854
rect 666 15850 807 15854
rect 841 15850 1026 15884
rect 666 15820 1026 15850
rect 603 15812 1026 15820
rect 603 15786 807 15812
rect 603 15752 632 15786
rect 666 15778 807 15786
rect 841 15778 1026 15812
rect 666 15752 1026 15778
rect 603 15740 1026 15752
rect 603 15718 807 15740
rect 603 15684 632 15718
rect 666 15706 807 15718
rect 841 15706 1026 15740
rect 666 15684 1026 15706
rect 603 15668 1026 15684
rect 603 15650 807 15668
rect 603 15616 632 15650
rect 666 15634 807 15650
rect 841 15634 1026 15668
rect 666 15616 1026 15634
rect 603 15596 1026 15616
rect 603 15582 807 15596
rect 603 15548 632 15582
rect 666 15562 807 15582
rect 841 15562 1026 15596
rect 666 15548 1026 15562
rect 603 15524 1026 15548
rect 603 15514 807 15524
rect 603 15480 632 15514
rect 666 15490 807 15514
rect 841 15490 1026 15524
rect 666 15480 1026 15490
rect 603 15452 1026 15480
rect 603 15446 807 15452
rect 603 15412 632 15446
rect 666 15418 807 15446
rect 841 15418 1026 15452
rect 666 15412 1026 15418
rect 603 15380 1026 15412
rect 603 15378 807 15380
rect 603 15344 632 15378
rect 666 15346 807 15378
rect 841 15346 1026 15380
rect 666 15344 1026 15346
rect 603 15310 1026 15344
rect 603 15276 632 15310
rect 666 15308 1026 15310
rect 666 15276 807 15308
rect 603 15274 807 15276
rect 841 15274 1026 15308
rect 603 15242 1026 15274
rect 603 15208 632 15242
rect 666 15236 1026 15242
rect 666 15208 807 15236
rect 603 15202 807 15208
rect 841 15202 1026 15236
rect 603 15174 1026 15202
rect 1119 34679 13887 34721
rect 1119 34645 1301 34679
rect 1339 34645 1373 34679
rect 1407 34645 1441 34679
rect 1479 34645 1509 34679
rect 1551 34645 1577 34679
rect 1623 34645 1645 34679
rect 1695 34645 1713 34679
rect 1767 34645 1781 34679
rect 1839 34645 1849 34679
rect 1911 34645 1917 34679
rect 1983 34645 1985 34679
rect 2019 34645 2021 34679
rect 2087 34645 2093 34679
rect 2155 34645 2165 34679
rect 2223 34645 2237 34679
rect 2291 34645 2309 34679
rect 2359 34645 2381 34679
rect 2427 34645 2453 34679
rect 2495 34645 2525 34679
rect 2563 34645 2597 34679
rect 2631 34645 2665 34679
rect 2703 34645 2733 34679
rect 2775 34645 2801 34679
rect 2847 34645 2869 34679
rect 2919 34645 2937 34679
rect 2991 34645 3005 34679
rect 3063 34645 3073 34679
rect 3135 34645 3141 34679
rect 3207 34645 3209 34679
rect 3243 34645 3245 34679
rect 3311 34645 3317 34679
rect 3379 34645 3389 34679
rect 3447 34645 3461 34679
rect 3515 34645 3533 34679
rect 3583 34645 3605 34679
rect 3651 34645 3677 34679
rect 3719 34645 3749 34679
rect 3787 34645 3821 34679
rect 3855 34645 3889 34679
rect 3927 34645 3957 34679
rect 3999 34645 4025 34679
rect 4071 34645 4093 34679
rect 4143 34645 4161 34679
rect 4215 34645 4229 34679
rect 4287 34645 4297 34679
rect 4359 34645 4365 34679
rect 4431 34645 4433 34679
rect 4467 34645 4469 34679
rect 4535 34645 4541 34679
rect 4603 34645 4613 34679
rect 4671 34645 4685 34679
rect 4739 34645 4757 34679
rect 4807 34645 4829 34679
rect 4875 34645 4901 34679
rect 4943 34645 4973 34679
rect 5011 34645 5045 34679
rect 5079 34645 5113 34679
rect 5151 34645 5181 34679
rect 5223 34645 5249 34679
rect 5295 34645 5317 34679
rect 5367 34645 5385 34679
rect 5439 34645 5453 34679
rect 5511 34645 5521 34679
rect 5583 34645 5589 34679
rect 5655 34645 5657 34679
rect 5691 34645 5693 34679
rect 5759 34645 5765 34679
rect 5827 34645 5837 34679
rect 5895 34645 5909 34679
rect 5963 34645 5981 34679
rect 6031 34645 6053 34679
rect 6099 34645 6125 34679
rect 6167 34645 6197 34679
rect 6235 34645 6269 34679
rect 6303 34645 6337 34679
rect 6375 34645 6405 34679
rect 6447 34645 6473 34679
rect 6519 34645 6541 34679
rect 6591 34645 6609 34679
rect 6663 34645 6677 34679
rect 6735 34645 6745 34679
rect 6807 34645 6813 34679
rect 6879 34645 6881 34679
rect 6915 34645 6917 34679
rect 6983 34645 6989 34679
rect 7051 34645 7061 34679
rect 7119 34645 7133 34679
rect 7187 34645 7205 34679
rect 7255 34645 7277 34679
rect 7323 34645 7349 34679
rect 7391 34645 7421 34679
rect 7459 34645 7493 34679
rect 7527 34645 7561 34679
rect 7599 34645 7629 34679
rect 7671 34645 7697 34679
rect 7743 34645 7765 34679
rect 7815 34645 7833 34679
rect 7887 34645 7901 34679
rect 7959 34645 7969 34679
rect 8031 34645 8037 34679
rect 8103 34645 8105 34679
rect 8139 34645 8141 34679
rect 8207 34645 8213 34679
rect 8275 34645 8285 34679
rect 8343 34645 8357 34679
rect 8411 34645 8429 34679
rect 8479 34645 8501 34679
rect 8547 34645 8573 34679
rect 8615 34645 8645 34679
rect 8683 34645 8717 34679
rect 8751 34645 8785 34679
rect 8823 34645 8853 34679
rect 8895 34645 8921 34679
rect 8967 34645 8989 34679
rect 9039 34645 9057 34679
rect 9111 34645 9125 34679
rect 9183 34645 9193 34679
rect 9255 34645 9261 34679
rect 9327 34645 9329 34679
rect 9363 34645 9365 34679
rect 9431 34645 9437 34679
rect 9499 34645 9509 34679
rect 9567 34645 9581 34679
rect 9635 34645 9653 34679
rect 9703 34645 9725 34679
rect 9771 34645 9797 34679
rect 9839 34645 9869 34679
rect 9907 34645 9941 34679
rect 9975 34645 10009 34679
rect 10047 34645 10077 34679
rect 10119 34645 10145 34679
rect 10191 34645 10213 34679
rect 10263 34645 10281 34679
rect 10335 34645 10349 34679
rect 10407 34645 10417 34679
rect 10479 34645 10485 34679
rect 10551 34645 10553 34679
rect 10587 34645 10589 34679
rect 10655 34645 10661 34679
rect 10723 34645 10733 34679
rect 10791 34645 10805 34679
rect 10859 34645 10877 34679
rect 10927 34645 10949 34679
rect 10995 34645 11021 34679
rect 11063 34645 11093 34679
rect 11131 34645 11165 34679
rect 11199 34645 11233 34679
rect 11271 34645 11301 34679
rect 11343 34645 11369 34679
rect 11415 34645 11437 34679
rect 11487 34645 11505 34679
rect 11559 34645 11573 34679
rect 11631 34645 11641 34679
rect 11703 34645 11709 34679
rect 11775 34645 11777 34679
rect 11811 34645 11813 34679
rect 11879 34645 11885 34679
rect 11947 34645 11957 34679
rect 12015 34645 12029 34679
rect 12083 34645 12101 34679
rect 12151 34645 12173 34679
rect 12219 34645 12245 34679
rect 12287 34645 12317 34679
rect 12355 34645 12389 34679
rect 12423 34645 12457 34679
rect 12495 34645 12525 34679
rect 12567 34645 12593 34679
rect 12639 34645 12661 34679
rect 12711 34645 12729 34679
rect 12783 34645 12797 34679
rect 12855 34645 12865 34679
rect 12927 34645 12933 34679
rect 12999 34645 13001 34679
rect 13035 34645 13037 34679
rect 13103 34645 13109 34679
rect 13171 34645 13181 34679
rect 13239 34645 13253 34679
rect 13307 34645 13325 34679
rect 13375 34645 13397 34679
rect 13443 34645 13469 34679
rect 13511 34645 13541 34679
rect 13579 34645 13613 34679
rect 13647 34645 13681 34679
rect 13719 34645 13887 34679
rect 1119 34603 13887 34645
rect 1119 34482 1237 34603
rect 1119 34428 1161 34482
rect 1195 34428 1237 34482
rect 1119 34410 1237 34428
rect 1119 34360 1161 34410
rect 1195 34360 1237 34410
rect 1119 34338 1237 34360
rect 1119 34292 1161 34338
rect 1195 34292 1237 34338
rect 1119 34266 1237 34292
rect 1119 34224 1161 34266
rect 1195 34224 1237 34266
rect 1119 34194 1237 34224
rect 1119 34156 1161 34194
rect 1195 34156 1237 34194
rect 1119 34122 1237 34156
rect 1119 34088 1161 34122
rect 1195 34088 1237 34122
rect 1119 34054 1237 34088
rect 1119 34016 1161 34054
rect 1195 34016 1237 34054
rect 1119 33986 1237 34016
rect 1119 33944 1161 33986
rect 1195 33944 1237 33986
rect 1119 33918 1237 33944
rect 1119 33872 1161 33918
rect 1195 33872 1237 33918
rect 1119 33850 1237 33872
rect 1119 33800 1161 33850
rect 1195 33800 1237 33850
rect 1119 33782 1237 33800
rect 1119 33728 1161 33782
rect 1195 33728 1237 33782
rect 1119 33714 1237 33728
rect 1119 33656 1161 33714
rect 1195 33656 1237 33714
rect 1119 33646 1237 33656
rect 1119 33584 1161 33646
rect 1195 33584 1237 33646
rect 1119 33578 1237 33584
rect 1119 33512 1161 33578
rect 1195 33512 1237 33578
rect 1119 33510 1237 33512
rect 1119 33476 1161 33510
rect 1195 33476 1237 33510
rect 1119 33474 1237 33476
rect 1119 33408 1161 33474
rect 1195 33408 1237 33474
rect 1119 33402 1237 33408
rect 1119 33340 1161 33402
rect 1195 33340 1237 33402
rect 1119 33330 1237 33340
rect 1119 33272 1161 33330
rect 1195 33272 1237 33330
rect 1119 33258 1237 33272
rect 1119 33204 1161 33258
rect 1195 33204 1237 33258
rect 1119 33186 1237 33204
rect 1119 33136 1161 33186
rect 1195 33136 1237 33186
rect 1119 33114 1237 33136
rect 1119 33068 1161 33114
rect 1195 33068 1237 33114
rect 1119 33042 1237 33068
rect 1119 33000 1161 33042
rect 1195 33000 1237 33042
rect 1119 32970 1237 33000
rect 1119 32932 1161 32970
rect 1195 32932 1237 32970
rect 1119 32898 1237 32932
rect 1119 32864 1161 32898
rect 1195 32864 1237 32898
rect 1119 32830 1237 32864
rect 1119 32792 1161 32830
rect 1195 32792 1237 32830
rect 1119 32762 1237 32792
rect 1119 32720 1161 32762
rect 1195 32720 1237 32762
rect 1119 32694 1237 32720
rect 1119 32648 1161 32694
rect 1195 32648 1237 32694
rect 1119 32626 1237 32648
rect 1119 32576 1161 32626
rect 1195 32576 1237 32626
rect 1119 32558 1237 32576
rect 1119 32504 1161 32558
rect 1195 32504 1237 32558
rect 1119 32490 1237 32504
rect 1119 32432 1161 32490
rect 1195 32432 1237 32490
rect 1119 32422 1237 32432
rect 1119 32360 1161 32422
rect 1195 32360 1237 32422
rect 1119 32354 1237 32360
rect 1119 32288 1161 32354
rect 1195 32288 1237 32354
rect 1119 32286 1237 32288
rect 1119 32252 1161 32286
rect 1195 32252 1237 32286
rect 1119 32250 1237 32252
rect 1119 32184 1161 32250
rect 1195 32184 1237 32250
rect 1119 32178 1237 32184
rect 1119 32116 1161 32178
rect 1195 32116 1237 32178
rect 1119 32106 1237 32116
rect 1119 32048 1161 32106
rect 1195 32048 1237 32106
rect 1119 32034 1237 32048
rect 1119 31980 1161 32034
rect 1195 31980 1237 32034
rect 1119 31962 1237 31980
rect 1119 31912 1161 31962
rect 1195 31912 1237 31962
rect 1119 31890 1237 31912
rect 1119 31844 1161 31890
rect 1195 31844 1237 31890
rect 1119 31818 1237 31844
rect 1119 31776 1161 31818
rect 1195 31776 1237 31818
rect 1119 31746 1237 31776
rect 1119 31708 1161 31746
rect 1195 31708 1237 31746
rect 1119 31674 1237 31708
rect 1119 31640 1161 31674
rect 1195 31640 1237 31674
rect 1119 31606 1237 31640
rect 1119 31568 1161 31606
rect 1195 31568 1237 31606
rect 1119 31538 1237 31568
rect 1119 31496 1161 31538
rect 1195 31496 1237 31538
rect 1119 31470 1237 31496
rect 1119 31424 1161 31470
rect 1195 31424 1237 31470
rect 1119 31402 1237 31424
rect 1119 31352 1161 31402
rect 1195 31352 1237 31402
rect 1119 31334 1237 31352
rect 1119 31280 1161 31334
rect 1195 31280 1237 31334
rect 1119 31266 1237 31280
rect 1119 31208 1161 31266
rect 1195 31208 1237 31266
rect 1119 31198 1237 31208
rect 1119 31136 1161 31198
rect 1195 31136 1237 31198
rect 1119 31130 1237 31136
rect 1119 31064 1161 31130
rect 1195 31064 1237 31130
rect 1119 31062 1237 31064
rect 1119 31028 1161 31062
rect 1195 31028 1237 31062
rect 1119 31026 1237 31028
rect 1119 30960 1161 31026
rect 1195 30960 1237 31026
rect 1119 30954 1237 30960
rect 1119 30892 1161 30954
rect 1195 30892 1237 30954
rect 1119 30882 1237 30892
rect 1119 30824 1161 30882
rect 1195 30824 1237 30882
rect 1119 30810 1237 30824
rect 1119 30756 1161 30810
rect 1195 30756 1237 30810
rect 1119 30738 1237 30756
rect 1119 30688 1161 30738
rect 1195 30688 1237 30738
rect 1119 30666 1237 30688
rect 1119 30620 1161 30666
rect 1195 30620 1237 30666
rect 1119 30594 1237 30620
rect 1119 30552 1161 30594
rect 1195 30552 1237 30594
rect 1119 30522 1237 30552
rect 1119 30484 1161 30522
rect 1195 30484 1237 30522
rect 1119 30450 1237 30484
rect 1119 30416 1161 30450
rect 1195 30416 1237 30450
rect 1119 30382 1237 30416
rect 1119 30344 1161 30382
rect 1195 30344 1237 30382
rect 1119 30314 1237 30344
rect 1119 30272 1161 30314
rect 1195 30272 1237 30314
rect 1119 30246 1237 30272
rect 1119 30200 1161 30246
rect 1195 30200 1237 30246
rect 1119 30178 1237 30200
rect 1119 30128 1161 30178
rect 1195 30128 1237 30178
rect 1119 30110 1237 30128
rect 1119 30056 1161 30110
rect 1195 30056 1237 30110
rect 1119 30042 1237 30056
rect 1119 29984 1161 30042
rect 1195 29984 1237 30042
rect 1119 29974 1237 29984
rect 1119 29912 1161 29974
rect 1195 29912 1237 29974
rect 1119 29906 1237 29912
rect 1119 29840 1161 29906
rect 1195 29840 1237 29906
rect 1119 29838 1237 29840
rect 1119 29804 1161 29838
rect 1195 29804 1237 29838
rect 1119 29802 1237 29804
rect 1119 29736 1161 29802
rect 1195 29736 1237 29802
rect 1119 29730 1237 29736
rect 1119 29668 1161 29730
rect 1195 29668 1237 29730
rect 1119 29658 1237 29668
rect 1119 29600 1161 29658
rect 1195 29600 1237 29658
rect 1119 29586 1237 29600
rect 1119 29532 1161 29586
rect 1195 29532 1237 29586
rect 1119 29514 1237 29532
rect 1119 29464 1161 29514
rect 1195 29464 1237 29514
rect 1119 29442 1237 29464
rect 1119 29396 1161 29442
rect 1195 29396 1237 29442
rect 1119 29370 1237 29396
rect 1119 29328 1161 29370
rect 1195 29328 1237 29370
rect 1119 29298 1237 29328
rect 1119 29260 1161 29298
rect 1195 29260 1237 29298
rect 1119 29226 1237 29260
rect 1119 29192 1161 29226
rect 1195 29192 1237 29226
rect 1119 29158 1237 29192
rect 1119 29120 1161 29158
rect 1195 29120 1237 29158
rect 1119 29090 1237 29120
rect 1119 29048 1161 29090
rect 1195 29048 1237 29090
rect 1119 29022 1237 29048
rect 1119 28976 1161 29022
rect 1195 28976 1237 29022
rect 1119 28954 1237 28976
rect 1119 28904 1161 28954
rect 1195 28904 1237 28954
rect 13769 34474 13887 34603
rect 13769 34423 13809 34474
rect 13843 34423 13887 34474
rect 13769 34402 13887 34423
rect 13769 34355 13809 34402
rect 13843 34355 13887 34402
rect 13769 34330 13887 34355
rect 13769 34287 13809 34330
rect 13843 34287 13887 34330
rect 13769 34258 13887 34287
rect 13769 34219 13809 34258
rect 13843 34219 13887 34258
rect 13769 34186 13887 34219
rect 13769 34151 13809 34186
rect 13843 34151 13887 34186
rect 13769 34117 13887 34151
rect 13769 34080 13809 34117
rect 13843 34080 13887 34117
rect 13769 34049 13887 34080
rect 13769 34008 13809 34049
rect 13843 34008 13887 34049
rect 13769 33981 13887 34008
rect 13769 33936 13809 33981
rect 13843 33936 13887 33981
rect 13769 33913 13887 33936
rect 13769 33864 13809 33913
rect 13843 33864 13887 33913
rect 13769 33845 13887 33864
rect 13769 33792 13809 33845
rect 13843 33792 13887 33845
rect 13769 33777 13887 33792
rect 13769 33720 13809 33777
rect 13843 33720 13887 33777
rect 13769 33709 13887 33720
rect 13769 33648 13809 33709
rect 13843 33648 13887 33709
rect 13769 33641 13887 33648
rect 13769 33576 13809 33641
rect 13843 33576 13887 33641
rect 13769 33573 13887 33576
rect 13769 33539 13809 33573
rect 13843 33539 13887 33573
rect 13769 33538 13887 33539
rect 13769 33471 13809 33538
rect 13843 33471 13887 33538
rect 13769 33466 13887 33471
rect 13769 33403 13809 33466
rect 13843 33403 13887 33466
rect 13769 33394 13887 33403
rect 13769 33335 13809 33394
rect 13843 33335 13887 33394
rect 13769 33322 13887 33335
rect 13769 33267 13809 33322
rect 13843 33267 13887 33322
rect 13769 33250 13887 33267
rect 13769 33199 13809 33250
rect 13843 33199 13887 33250
rect 13769 33178 13887 33199
rect 13769 33131 13809 33178
rect 13843 33131 13887 33178
rect 13769 33106 13887 33131
rect 13769 33063 13809 33106
rect 13843 33063 13887 33106
rect 13769 33034 13887 33063
rect 13769 32995 13809 33034
rect 13843 32995 13887 33034
rect 13769 32962 13887 32995
rect 13769 32927 13809 32962
rect 13843 32927 13887 32962
rect 13769 32893 13887 32927
rect 13769 32856 13809 32893
rect 13843 32856 13887 32893
rect 13769 32825 13887 32856
rect 13769 32784 13809 32825
rect 13843 32784 13887 32825
rect 13769 32757 13887 32784
rect 13769 32712 13809 32757
rect 13843 32712 13887 32757
rect 13769 32689 13887 32712
rect 13769 32640 13809 32689
rect 13843 32640 13887 32689
rect 13769 32621 13887 32640
rect 13769 32568 13809 32621
rect 13843 32568 13887 32621
rect 13769 32553 13887 32568
rect 13769 32496 13809 32553
rect 13843 32496 13887 32553
rect 13769 32485 13887 32496
rect 13769 32424 13809 32485
rect 13843 32424 13887 32485
rect 13769 32417 13887 32424
rect 13769 32352 13809 32417
rect 13843 32352 13887 32417
rect 13769 32349 13887 32352
rect 13769 32315 13809 32349
rect 13843 32315 13887 32349
rect 13769 32314 13887 32315
rect 13769 32247 13809 32314
rect 13843 32247 13887 32314
rect 13769 32242 13887 32247
rect 13769 32179 13809 32242
rect 13843 32179 13887 32242
rect 13769 32170 13887 32179
rect 13769 32111 13809 32170
rect 13843 32111 13887 32170
rect 13769 32098 13887 32111
rect 13769 32043 13809 32098
rect 13843 32043 13887 32098
rect 13769 32026 13887 32043
rect 13769 31975 13809 32026
rect 13843 31975 13887 32026
rect 13769 31954 13887 31975
rect 13769 31907 13809 31954
rect 13843 31907 13887 31954
rect 13769 31882 13887 31907
rect 13769 31839 13809 31882
rect 13843 31839 13887 31882
rect 13769 31810 13887 31839
rect 13769 31771 13809 31810
rect 13843 31771 13887 31810
rect 13769 31738 13887 31771
rect 13769 31703 13809 31738
rect 13843 31703 13887 31738
rect 13769 31669 13887 31703
rect 13769 31632 13809 31669
rect 13843 31632 13887 31669
rect 13769 31601 13887 31632
rect 13769 31560 13809 31601
rect 13843 31560 13887 31601
rect 13769 31533 13887 31560
rect 13769 31488 13809 31533
rect 13843 31488 13887 31533
rect 13769 31465 13887 31488
rect 13769 31416 13809 31465
rect 13843 31416 13887 31465
rect 13769 31397 13887 31416
rect 13769 31344 13809 31397
rect 13843 31344 13887 31397
rect 13769 31329 13887 31344
rect 13769 31272 13809 31329
rect 13843 31272 13887 31329
rect 13769 31261 13887 31272
rect 13769 31200 13809 31261
rect 13843 31200 13887 31261
rect 13769 31193 13887 31200
rect 13769 31128 13809 31193
rect 13843 31128 13887 31193
rect 13769 31125 13887 31128
rect 13769 31091 13809 31125
rect 13843 31091 13887 31125
rect 13769 31090 13887 31091
rect 13769 31023 13809 31090
rect 13843 31023 13887 31090
rect 13769 31018 13887 31023
rect 13769 30955 13809 31018
rect 13843 30955 13887 31018
rect 13769 30946 13887 30955
rect 13769 30887 13809 30946
rect 13843 30887 13887 30946
rect 13769 30874 13887 30887
rect 13769 30819 13809 30874
rect 13843 30819 13887 30874
rect 13769 30802 13887 30819
rect 13769 30751 13809 30802
rect 13843 30751 13887 30802
rect 13769 30730 13887 30751
rect 13769 30683 13809 30730
rect 13843 30683 13887 30730
rect 13769 30658 13887 30683
rect 13769 30615 13809 30658
rect 13843 30615 13887 30658
rect 13769 30586 13887 30615
rect 13769 30547 13809 30586
rect 13843 30547 13887 30586
rect 13769 30514 13887 30547
rect 13769 30479 13809 30514
rect 13843 30479 13887 30514
rect 13769 30445 13887 30479
rect 13769 30408 13809 30445
rect 13843 30408 13887 30445
rect 13769 30377 13887 30408
rect 13769 30336 13809 30377
rect 13843 30336 13887 30377
rect 13769 30309 13887 30336
rect 13769 30264 13809 30309
rect 13843 30264 13887 30309
rect 13769 30241 13887 30264
rect 13769 30192 13809 30241
rect 13843 30192 13887 30241
rect 13769 30173 13887 30192
rect 13769 30120 13809 30173
rect 13843 30120 13887 30173
rect 13769 30105 13887 30120
rect 13769 30048 13809 30105
rect 13843 30048 13887 30105
rect 13769 30037 13887 30048
rect 13769 29976 13809 30037
rect 13843 29976 13887 30037
rect 13769 29969 13887 29976
rect 13769 29904 13809 29969
rect 13843 29904 13887 29969
rect 13769 29901 13887 29904
rect 13769 29867 13809 29901
rect 13843 29867 13887 29901
rect 13769 29866 13887 29867
rect 13769 29799 13809 29866
rect 13843 29799 13887 29866
rect 13769 29794 13887 29799
rect 13769 29731 13809 29794
rect 13843 29731 13887 29794
rect 13769 29722 13887 29731
rect 13769 29663 13809 29722
rect 13843 29663 13887 29722
rect 13769 29650 13887 29663
rect 13769 29595 13809 29650
rect 13843 29595 13887 29650
rect 13769 29578 13887 29595
rect 13769 29527 13809 29578
rect 13843 29527 13887 29578
rect 13769 29506 13887 29527
rect 13769 29459 13809 29506
rect 13843 29459 13887 29506
rect 13769 29434 13887 29459
rect 13769 29391 13809 29434
rect 13843 29391 13887 29434
rect 13769 29362 13887 29391
rect 13769 29323 13809 29362
rect 13843 29323 13887 29362
rect 13769 29290 13887 29323
rect 13769 29255 13809 29290
rect 13843 29255 13887 29290
rect 13769 29221 13887 29255
rect 13769 29184 13809 29221
rect 13843 29184 13887 29221
rect 13769 29153 13887 29184
rect 13769 29112 13809 29153
rect 13843 29112 13887 29153
rect 13769 29085 13887 29112
rect 13769 29040 13809 29085
rect 13843 29040 13887 29085
rect 13769 29017 13887 29040
rect 13769 28968 13809 29017
rect 13843 28968 13887 29017
rect 13769 28949 13887 28968
rect 1119 28886 1237 28904
rect 1119 28832 1161 28886
rect 1195 28832 1237 28886
rect 1119 28818 1237 28832
rect 1119 28760 1161 28818
rect 1195 28760 1237 28818
rect 1119 28750 1237 28760
rect 1119 28688 1161 28750
rect 1195 28688 1237 28750
rect 1119 28682 1237 28688
rect 1119 28616 1161 28682
rect 1195 28616 1237 28682
rect 1119 28614 1237 28616
rect 1119 28580 1161 28614
rect 1195 28580 1237 28614
rect 1119 28578 1237 28580
rect 1119 28512 1161 28578
rect 1195 28512 1237 28578
rect 1119 28506 1237 28512
rect 1119 28444 1161 28506
rect 1195 28444 1237 28506
rect 1119 28434 1237 28444
rect 1119 28376 1161 28434
rect 1195 28376 1237 28434
rect 1119 28362 1237 28376
rect 1119 28308 1161 28362
rect 1195 28308 1237 28362
rect 1119 28290 1237 28308
rect 1119 28240 1161 28290
rect 1195 28240 1237 28290
rect 1119 28218 1237 28240
rect 1119 28172 1161 28218
rect 1195 28172 1237 28218
rect 1119 28146 1237 28172
rect 1119 28104 1161 28146
rect 1195 28104 1237 28146
rect 1119 28074 1237 28104
rect 1119 28036 1161 28074
rect 1195 28036 1237 28074
rect 1119 28002 1237 28036
rect 1119 27968 1161 28002
rect 1195 27968 1237 28002
rect 1119 27934 1237 27968
rect 1119 27896 1161 27934
rect 1195 27896 1237 27934
rect 1119 27866 1237 27896
rect 1119 27824 1161 27866
rect 1195 27824 1237 27866
rect 1119 27798 1237 27824
rect 1119 27752 1161 27798
rect 1195 27752 1237 27798
rect 1119 27730 1237 27752
rect 1119 27680 1161 27730
rect 1195 27680 1237 27730
rect 1119 27662 1237 27680
rect 1119 27608 1161 27662
rect 1195 27608 1237 27662
rect 1119 27594 1237 27608
rect 1119 27536 1161 27594
rect 1195 27536 1237 27594
rect 1119 27526 1237 27536
rect 1119 27464 1161 27526
rect 1195 27464 1237 27526
rect 1119 27458 1237 27464
rect 1119 27392 1161 27458
rect 1195 27392 1237 27458
rect 1119 27390 1237 27392
rect 1119 27356 1161 27390
rect 1195 27356 1237 27390
rect 1119 27354 1237 27356
rect 1119 27288 1161 27354
rect 1195 27288 1237 27354
rect 1119 27282 1237 27288
rect 1119 27220 1161 27282
rect 1195 27220 1237 27282
rect 1119 27210 1237 27220
rect 1119 27152 1161 27210
rect 1195 27152 1237 27210
rect 1119 27138 1237 27152
rect 1119 27084 1161 27138
rect 1195 27084 1237 27138
rect 1119 27066 1237 27084
rect 1119 27016 1161 27066
rect 1195 27016 1237 27066
rect 1659 28879 13357 28909
rect 1659 28875 2119 28879
rect 12897 28875 13357 28879
rect 1659 28553 1982 28875
rect 13032 28553 13357 28875
rect 1659 28505 2119 28553
rect 12897 28505 13357 28553
rect 1659 28489 13357 28505
rect 1659 28422 1726 28489
rect 1976 28482 13357 28489
rect 1976 28475 13031 28482
rect 1976 28422 2093 28475
rect 1659 27504 1689 28422
rect 2063 27504 2093 28422
rect 12923 28422 13031 28475
rect 13281 28422 13357 28482
rect 2156 28172 12840 28368
rect 2156 27758 2382 28172
rect 12614 27758 12840 28172
rect 2156 27556 12840 27758
rect 1659 27447 1726 27504
rect 1976 27451 2093 27504
rect 12923 27504 12953 28422
rect 13327 27504 13357 28422
rect 12923 27451 13031 27504
rect 1976 27447 13031 27451
rect 1659 27440 13031 27447
rect 13281 27440 13357 27504
rect 1659 27421 13357 27440
rect 1659 27334 2119 27421
rect 12897 27334 13357 27421
rect 1659 27084 1985 27334
rect 13035 27084 13357 27334
rect 1659 27047 2119 27084
rect 12897 27047 13357 27084
rect 1659 27017 13357 27047
rect 13769 28896 13809 28949
rect 13843 28896 13887 28949
rect 13769 28881 13887 28896
rect 13769 28824 13809 28881
rect 13843 28824 13887 28881
rect 13769 28813 13887 28824
rect 13769 28752 13809 28813
rect 13843 28752 13887 28813
rect 13769 28745 13887 28752
rect 13769 28711 13809 28745
rect 13843 28711 13887 28745
rect 13769 28677 13887 28711
rect 13769 28643 13809 28677
rect 13843 28643 13887 28677
rect 13769 28609 13887 28643
rect 13769 28575 13809 28609
rect 13843 28575 13887 28609
rect 13769 28541 13887 28575
rect 13769 28507 13809 28541
rect 13843 28507 13887 28541
rect 13769 28473 13887 28507
rect 13769 28439 13809 28473
rect 13843 28439 13887 28473
rect 13769 28405 13887 28439
rect 13769 28371 13809 28405
rect 13843 28371 13887 28405
rect 13769 28337 13887 28371
rect 13769 28303 13809 28337
rect 13843 28303 13887 28337
rect 13769 28269 13887 28303
rect 13769 28235 13809 28269
rect 13843 28235 13887 28269
rect 13769 28201 13887 28235
rect 13769 28167 13809 28201
rect 13843 28167 13887 28201
rect 13769 28133 13887 28167
rect 13769 28099 13809 28133
rect 13843 28099 13887 28133
rect 13769 28065 13887 28099
rect 13769 28031 13809 28065
rect 13843 28031 13887 28065
rect 13769 27997 13887 28031
rect 13769 27963 13809 27997
rect 13843 27963 13887 27997
rect 13769 27929 13887 27963
rect 13769 27895 13809 27929
rect 13843 27895 13887 27929
rect 13769 27861 13887 27895
rect 13769 27827 13809 27861
rect 13843 27827 13887 27861
rect 13769 27793 13887 27827
rect 13769 27759 13809 27793
rect 13843 27759 13887 27793
rect 13769 27725 13887 27759
rect 13769 27691 13809 27725
rect 13843 27691 13887 27725
rect 13769 27657 13887 27691
rect 13769 27623 13809 27657
rect 13843 27623 13887 27657
rect 13769 27589 13887 27623
rect 13769 27555 13809 27589
rect 13843 27555 13887 27589
rect 13769 27521 13887 27555
rect 13769 27487 13809 27521
rect 13843 27487 13887 27521
rect 13769 27453 13887 27487
rect 13769 27419 13809 27453
rect 13843 27419 13887 27453
rect 13769 27385 13887 27419
rect 13769 27351 13809 27385
rect 13843 27351 13887 27385
rect 13769 27317 13887 27351
rect 13769 27283 13809 27317
rect 13843 27283 13887 27317
rect 13769 27249 13887 27283
rect 13769 27215 13809 27249
rect 13843 27215 13887 27249
rect 13769 27181 13887 27215
rect 13769 27147 13809 27181
rect 13843 27147 13887 27181
rect 13769 27113 13887 27147
rect 13769 27079 13809 27113
rect 13843 27079 13887 27113
rect 13769 27045 13887 27079
rect 1119 26994 1237 27016
rect 1119 26948 1161 26994
rect 1195 26948 1237 26994
rect 1119 26922 1237 26948
rect 1119 26880 1161 26922
rect 1195 26880 1237 26922
rect 1119 26850 1237 26880
rect 1119 26812 1161 26850
rect 1195 26812 1237 26850
rect 1119 26778 1237 26812
rect 1119 26744 1161 26778
rect 1195 26744 1237 26778
rect 1119 26710 1237 26744
rect 1119 26672 1161 26710
rect 1195 26672 1237 26710
rect 1119 26642 1237 26672
rect 1119 26600 1161 26642
rect 1195 26600 1237 26642
rect 13769 27011 13809 27045
rect 13843 27011 13887 27045
rect 13769 26977 13887 27011
rect 13769 26943 13809 26977
rect 13843 26943 13887 26977
rect 13769 26909 13887 26943
rect 13769 26875 13809 26909
rect 13843 26875 13887 26909
rect 13769 26841 13887 26875
rect 13769 26807 13809 26841
rect 13843 26807 13887 26841
rect 13769 26773 13887 26807
rect 13769 26739 13809 26773
rect 13843 26739 13887 26773
rect 13769 26705 13887 26739
rect 13769 26671 13809 26705
rect 13843 26671 13887 26705
rect 13769 26637 13887 26671
rect 13769 26613 13809 26637
rect 1119 26574 1237 26600
rect 1119 26528 1161 26574
rect 1195 26528 1237 26574
rect 1119 26506 1237 26528
rect 1119 26456 1161 26506
rect 1195 26456 1237 26506
rect 1119 26438 1237 26456
rect 1119 26384 1161 26438
rect 1195 26384 1237 26438
rect 1119 26370 1237 26384
rect 1119 26312 1161 26370
rect 1195 26312 1237 26370
rect 1119 26302 1237 26312
rect 1119 26240 1161 26302
rect 1195 26240 1237 26302
rect 1119 26234 1237 26240
rect 1119 26168 1161 26234
rect 1195 26168 1237 26234
rect 1119 26166 1237 26168
rect 1119 26132 1161 26166
rect 1195 26132 1237 26166
rect 1119 26130 1237 26132
rect 1119 26064 1161 26130
rect 1195 26064 1237 26130
rect 1119 26058 1237 26064
rect 1119 25996 1161 26058
rect 1195 25996 1237 26058
rect 1119 25986 1237 25996
rect 1119 25928 1161 25986
rect 1195 25928 1237 25986
rect 1119 25914 1237 25928
rect 1119 25860 1161 25914
rect 1195 25860 1237 25914
rect 1119 25842 1237 25860
rect 1119 25792 1161 25842
rect 1195 25792 1237 25842
rect 1119 25770 1237 25792
rect 1119 25724 1161 25770
rect 1195 25724 1237 25770
rect 1119 25698 1237 25724
rect 1119 25656 1161 25698
rect 1195 25656 1237 25698
rect 1119 25626 1237 25656
rect 1119 25588 1161 25626
rect 1195 25588 1237 25626
rect 1119 25554 1237 25588
rect 1119 25520 1161 25554
rect 1195 25520 1237 25554
rect 1119 25486 1237 25520
rect 1119 25448 1161 25486
rect 1195 25448 1237 25486
rect 1119 25418 1237 25448
rect 1119 25376 1161 25418
rect 1195 25376 1237 25418
rect 1119 25350 1237 25376
rect 1119 25304 1161 25350
rect 1195 25304 1237 25350
rect 1119 25282 1237 25304
rect 1119 25232 1161 25282
rect 1195 25232 1237 25282
rect 1119 25214 1237 25232
rect 1119 25160 1161 25214
rect 1195 25160 1237 25214
rect 1119 25146 1237 25160
rect 1119 25088 1161 25146
rect 1195 25088 1237 25146
rect 1119 25078 1237 25088
rect 1119 25016 1161 25078
rect 1195 25016 1237 25078
rect 1119 25010 1237 25016
rect 1119 24944 1161 25010
rect 1195 24944 1237 25010
rect 1119 24942 1237 24944
rect 1119 24908 1161 24942
rect 1195 24908 1237 24942
rect 1119 24906 1237 24908
rect 1119 24840 1161 24906
rect 1195 24840 1237 24906
rect 1119 24834 1237 24840
rect 1119 24772 1161 24834
rect 1195 24772 1237 24834
rect 1698 26603 13809 26613
rect 13843 26603 13887 26637
rect 1698 26569 13887 26603
rect 1698 26535 13809 26569
rect 13843 26535 13887 26569
rect 1698 26501 13887 26535
rect 1698 26467 13809 26501
rect 13843 26467 13887 26501
rect 1698 26433 13887 26467
rect 1698 26399 13809 26433
rect 13843 26399 13887 26433
rect 1698 26365 13887 26399
rect 1698 26331 13809 26365
rect 13843 26331 13887 26365
rect 1698 26297 13887 26331
rect 1698 26263 13809 26297
rect 13843 26263 13887 26297
rect 1698 26229 13887 26263
rect 1698 26195 13809 26229
rect 13843 26195 13887 26229
rect 1698 26161 13887 26195
rect 1698 26127 13809 26161
rect 13843 26127 13887 26161
rect 1698 26093 13887 26127
rect 1698 26080 13809 26093
rect 1698 25313 2270 26080
rect 12712 26059 13809 26080
rect 13843 26059 13887 26093
rect 12712 26025 13887 26059
rect 12712 25991 13809 26025
rect 13843 25991 13887 26025
rect 12712 25957 13887 25991
rect 12712 25923 13809 25957
rect 13843 25923 13887 25957
rect 12712 25889 13887 25923
rect 12712 25855 13809 25889
rect 13843 25855 13887 25889
rect 12712 25821 13887 25855
rect 12712 25787 13809 25821
rect 13843 25787 13887 25821
rect 12712 25753 13887 25787
rect 12712 25719 13809 25753
rect 13843 25719 13887 25753
rect 12712 25685 13887 25719
rect 12712 25651 13809 25685
rect 13843 25651 13887 25685
rect 12712 25617 13887 25651
rect 12712 25583 13809 25617
rect 13843 25583 13887 25617
rect 12712 25549 13887 25583
rect 12712 25515 13809 25549
rect 13843 25515 13887 25549
rect 12712 25481 13887 25515
rect 12712 25447 13809 25481
rect 13843 25447 13887 25481
rect 12712 25413 13887 25447
rect 12712 25379 13809 25413
rect 13843 25379 13887 25413
rect 12712 25345 13887 25379
rect 12712 25313 13809 25345
rect 1698 25311 13809 25313
rect 13843 25311 13887 25345
rect 1698 25277 13887 25311
rect 1698 25243 13809 25277
rect 13843 25243 13887 25277
rect 1698 25209 13887 25243
rect 1698 25175 13809 25209
rect 13843 25175 13887 25209
rect 1698 25141 13887 25175
rect 1698 25107 13809 25141
rect 13843 25107 13887 25141
rect 1698 25073 13887 25107
rect 1698 25039 13809 25073
rect 13843 25039 13887 25073
rect 1698 25005 13887 25039
rect 1698 24971 13809 25005
rect 13843 24971 13887 25005
rect 1698 24937 13887 24971
rect 1698 24903 13809 24937
rect 13843 24903 13887 24937
rect 1698 24869 13887 24903
rect 1698 24835 13809 24869
rect 13843 24835 13887 24869
rect 1698 24801 13887 24835
rect 1698 24780 13809 24801
rect 1119 24762 1237 24772
rect 1119 24704 1161 24762
rect 1195 24704 1237 24762
rect 1119 24690 1237 24704
rect 1119 24636 1161 24690
rect 1195 24636 1237 24690
rect 1119 24618 1237 24636
rect 1119 24568 1161 24618
rect 1195 24568 1237 24618
rect 1119 24546 1237 24568
rect 1119 24500 1161 24546
rect 1195 24500 1237 24546
rect 1119 24474 1237 24500
rect 1119 24432 1161 24474
rect 1195 24432 1237 24474
rect 1119 24402 1237 24432
rect 1119 24364 1161 24402
rect 1195 24364 1237 24402
rect 1119 24330 1237 24364
rect 1119 24296 1161 24330
rect 1195 24296 1237 24330
rect 1119 24262 1237 24296
rect 1119 24224 1161 24262
rect 1195 24224 1237 24262
rect 1119 24194 1237 24224
rect 1119 24152 1161 24194
rect 1195 24152 1237 24194
rect 1119 24126 1237 24152
rect 1119 24080 1161 24126
rect 1195 24080 1237 24126
rect 1119 24058 1237 24080
rect 1119 24008 1161 24058
rect 1195 24008 1237 24058
rect 1119 23990 1237 24008
rect 1119 23936 1161 23990
rect 1195 23936 1237 23990
rect 1119 23922 1237 23936
rect 1119 23864 1161 23922
rect 1195 23864 1237 23922
rect 1119 23854 1237 23864
rect 1119 23792 1161 23854
rect 1195 23792 1237 23854
rect 1119 23786 1237 23792
rect 1119 23720 1161 23786
rect 1195 23720 1237 23786
rect 1119 23718 1237 23720
rect 1119 23684 1161 23718
rect 1195 23684 1237 23718
rect 1119 23682 1237 23684
rect 1119 23616 1161 23682
rect 1195 23616 1237 23682
rect 1119 23610 1237 23616
rect 1119 23548 1161 23610
rect 1195 23548 1237 23610
rect 1119 23538 1237 23548
rect 1119 23480 1161 23538
rect 1195 23480 1237 23538
rect 1119 23466 1237 23480
rect 1119 23412 1161 23466
rect 1195 23412 1237 23466
rect 1119 23394 1237 23412
rect 1119 23344 1161 23394
rect 1195 23344 1237 23394
rect 1119 23322 1237 23344
rect 1119 23276 1161 23322
rect 1195 23276 1237 23322
rect 1119 23250 1237 23276
rect 1119 23208 1161 23250
rect 1195 23208 1237 23250
rect 1119 23178 1237 23208
rect 1119 23140 1161 23178
rect 1195 23140 1237 23178
rect 1119 23106 1237 23140
rect 1119 23072 1161 23106
rect 1195 23072 1237 23106
rect 1119 23038 1237 23072
rect 1119 23000 1161 23038
rect 1195 23000 1237 23038
rect 1119 22970 1237 23000
rect 1119 22928 1161 22970
rect 1195 22928 1237 22970
rect 1119 22902 1237 22928
rect 1119 22856 1161 22902
rect 1195 22856 1237 22902
rect 1119 22834 1237 22856
rect 1119 22784 1161 22834
rect 1195 22784 1237 22834
rect 1119 22766 1237 22784
rect 1119 22712 1161 22766
rect 1195 22712 1237 22766
rect 1119 22698 1237 22712
rect 1119 22640 1161 22698
rect 1195 22640 1237 22698
rect 1119 22630 1237 22640
rect 1119 22568 1161 22630
rect 1195 22568 1237 22630
rect 1119 22562 1237 22568
rect 1119 22496 1161 22562
rect 1195 22496 1237 22562
rect 1119 22494 1237 22496
rect 1119 22460 1161 22494
rect 1195 22460 1237 22494
rect 1119 22458 1237 22460
rect 1119 22392 1161 22458
rect 1195 22392 1237 22458
rect 1119 22386 1237 22392
rect 1119 22324 1161 22386
rect 1195 22324 1237 22386
rect 1119 22314 1237 22324
rect 1119 22256 1161 22314
rect 1195 22256 1237 22314
rect 1119 22242 1237 22256
rect 1119 22188 1161 22242
rect 1195 22188 1237 22242
rect 1119 22170 1237 22188
rect 1119 22120 1161 22170
rect 1195 22120 1237 22170
rect 1119 22098 1237 22120
rect 1119 22052 1161 22098
rect 1195 22052 1237 22098
rect 1119 22026 1237 22052
rect 1119 21984 1161 22026
rect 1195 21984 1237 22026
rect 1119 21954 1237 21984
rect 1119 21916 1161 21954
rect 1195 21916 1237 21954
rect 1119 21882 1237 21916
rect 1119 21848 1161 21882
rect 1195 21848 1237 21882
rect 1119 21814 1237 21848
rect 1119 21776 1161 21814
rect 1195 21776 1237 21814
rect 1119 21746 1237 21776
rect 1119 21704 1161 21746
rect 1195 21704 1237 21746
rect 1119 21678 1237 21704
rect 1119 21632 1161 21678
rect 1195 21632 1237 21678
rect 1119 21610 1237 21632
rect 1119 21560 1161 21610
rect 1195 21560 1237 21610
rect 1119 21542 1237 21560
rect 1119 21488 1161 21542
rect 1195 21488 1237 21542
rect 1119 21474 1237 21488
rect 1119 21416 1161 21474
rect 1195 21416 1237 21474
rect 1119 21406 1237 21416
rect 1119 21344 1161 21406
rect 1195 21344 1237 21406
rect 1119 21338 1237 21344
rect 1119 21272 1161 21338
rect 1195 21272 1237 21338
rect 1119 21270 1237 21272
rect 1119 21236 1161 21270
rect 1195 21236 1237 21270
rect 1119 21234 1237 21236
rect 1119 21168 1161 21234
rect 1195 21168 1237 21234
rect 1119 21162 1237 21168
rect 1119 21100 1161 21162
rect 1195 21100 1237 21162
rect 1119 21090 1237 21100
rect 1119 21032 1161 21090
rect 1195 21032 1237 21090
rect 1119 21018 1237 21032
rect 1119 20964 1161 21018
rect 1195 20964 1237 21018
rect 1119 20946 1237 20964
rect 1119 20896 1161 20946
rect 1195 20896 1237 20946
rect 1119 20874 1237 20896
rect 1119 20828 1161 20874
rect 1195 20828 1237 20874
rect 1119 20802 1237 20828
rect 1119 20760 1161 20802
rect 1195 20760 1237 20802
rect 1119 20730 1237 20760
rect 1119 20692 1161 20730
rect 1195 20692 1237 20730
rect 1119 20658 1237 20692
rect 1119 20624 1161 20658
rect 1195 20624 1237 20658
rect 1119 20590 1237 20624
rect 1119 20552 1161 20590
rect 1195 20552 1237 20590
rect 1119 20522 1237 20552
rect 1119 20480 1161 20522
rect 1195 20480 1237 20522
rect 1119 20454 1237 20480
rect 1119 20408 1161 20454
rect 1195 20408 1237 20454
rect 1119 20386 1237 20408
rect 1119 20336 1161 20386
rect 1195 20336 1237 20386
rect 1119 20318 1237 20336
rect 1119 20264 1161 20318
rect 1195 20264 1237 20318
rect 1119 20250 1237 20264
rect 1119 20192 1161 20250
rect 1195 20192 1237 20250
rect 1119 20182 1237 20192
rect 1119 20120 1161 20182
rect 1195 20120 1237 20182
rect 1119 20114 1237 20120
rect 1119 20048 1161 20114
rect 1195 20048 1237 20114
rect 1119 20046 1237 20048
rect 1119 20012 1161 20046
rect 1195 20012 1237 20046
rect 1119 20010 1237 20012
rect 1119 19944 1161 20010
rect 1195 19944 1237 20010
rect 1119 19938 1237 19944
rect 1119 19876 1161 19938
rect 1195 19876 1237 19938
rect 1119 19866 1237 19876
rect 1119 19808 1161 19866
rect 1195 19808 1237 19866
rect 1119 19794 1237 19808
rect 1119 19740 1161 19794
rect 1195 19740 1237 19794
rect 1119 19722 1237 19740
rect 1119 19672 1161 19722
rect 1195 19672 1237 19722
rect 1119 19650 1237 19672
rect 1119 19604 1161 19650
rect 1195 19604 1237 19650
rect 1119 19578 1237 19604
rect 1119 19536 1161 19578
rect 1195 19536 1237 19578
rect 1119 19506 1237 19536
rect 1119 19468 1161 19506
rect 1195 19468 1237 19506
rect 1119 19434 1237 19468
rect 1119 19400 1161 19434
rect 1195 19400 1237 19434
rect 1119 19366 1237 19400
rect 1119 19328 1161 19366
rect 1195 19328 1237 19366
rect 1119 19298 1237 19328
rect 1119 19256 1161 19298
rect 1195 19256 1237 19298
rect 1119 19230 1237 19256
rect 1119 19184 1161 19230
rect 1195 19184 1237 19230
rect 1119 19162 1237 19184
rect 1119 19112 1161 19162
rect 1195 19112 1237 19162
rect 1119 19094 1237 19112
rect 1119 19040 1161 19094
rect 1195 19040 1237 19094
rect 1119 19026 1237 19040
rect 1119 18968 1161 19026
rect 1195 18968 1237 19026
rect 1119 18958 1237 18968
rect 1119 18896 1161 18958
rect 1195 18896 1237 18958
rect 1119 18890 1237 18896
rect 1119 18824 1161 18890
rect 1195 18824 1237 18890
rect 1119 18822 1237 18824
rect 1119 18788 1161 18822
rect 1195 18788 1237 18822
rect 1119 18786 1237 18788
rect 1119 18720 1161 18786
rect 1195 18720 1237 18786
rect 1119 18714 1237 18720
rect 1119 18652 1161 18714
rect 1195 18652 1237 18714
rect 1119 18642 1237 18652
rect 1119 18584 1161 18642
rect 1195 18584 1237 18642
rect 1119 18570 1237 18584
rect 1119 18516 1161 18570
rect 1195 18516 1237 18570
rect 1119 18498 1237 18516
rect 1119 18448 1161 18498
rect 1195 18448 1237 18498
rect 1119 18426 1237 18448
rect 1119 18380 1161 18426
rect 1195 18380 1237 18426
rect 1119 18354 1237 18380
rect 1119 18312 1161 18354
rect 1195 18312 1237 18354
rect 1119 18282 1237 18312
rect 1119 18244 1161 18282
rect 1195 18244 1237 18282
rect 1119 18210 1237 18244
rect 1119 18176 1161 18210
rect 1195 18176 1237 18210
rect 1119 18142 1237 18176
rect 1119 18104 1161 18142
rect 1195 18104 1237 18142
rect 1119 18074 1237 18104
rect 1119 18032 1161 18074
rect 1195 18032 1237 18074
rect 1119 18006 1237 18032
rect 1119 17960 1161 18006
rect 1195 17960 1237 18006
rect 1119 17938 1237 17960
rect 1119 17888 1161 17938
rect 1195 17888 1237 17938
rect 1119 17870 1237 17888
rect 1119 17816 1161 17870
rect 1195 17816 1237 17870
rect 1119 17802 1237 17816
rect 1119 17744 1161 17802
rect 1195 17744 1237 17802
rect 1119 17734 1237 17744
rect 1119 17672 1161 17734
rect 1195 17672 1237 17734
rect 1119 17666 1237 17672
rect 1119 17600 1161 17666
rect 1195 17600 1237 17666
rect 1119 17598 1237 17600
rect 1119 17564 1161 17598
rect 1195 17564 1237 17598
rect 1119 17562 1237 17564
rect 1119 17496 1161 17562
rect 1195 17496 1237 17562
rect 1119 17490 1237 17496
rect 1119 17428 1161 17490
rect 1195 17428 1237 17490
rect 1119 17418 1237 17428
rect 1119 17360 1161 17418
rect 1195 17360 1237 17418
rect 1119 17346 1237 17360
rect 1119 17292 1161 17346
rect 1195 17292 1237 17346
rect 1119 17274 1237 17292
rect 1119 17224 1161 17274
rect 1195 17224 1237 17274
rect 1119 17202 1237 17224
rect 1119 17156 1161 17202
rect 1195 17156 1237 17202
rect 1119 17130 1237 17156
rect 1119 17088 1161 17130
rect 1195 17088 1237 17130
rect 1119 17058 1237 17088
rect 1119 17020 1161 17058
rect 1195 17020 1237 17058
rect 1119 16986 1237 17020
rect 1119 16952 1161 16986
rect 1195 16952 1237 16986
rect 1119 16918 1237 16952
rect 1119 16880 1161 16918
rect 1195 16880 1237 16918
rect 1119 16850 1237 16880
rect 1119 16808 1161 16850
rect 1195 16808 1237 16850
rect 1119 16782 1237 16808
rect 1119 16736 1161 16782
rect 1195 16736 1237 16782
rect 1119 16714 1237 16736
rect 1119 16664 1161 16714
rect 1195 16664 1237 16714
rect 1119 16646 1237 16664
rect 1119 16592 1161 16646
rect 1195 16592 1237 16646
rect 1119 16578 1237 16592
rect 1119 16520 1161 16578
rect 1195 16520 1237 16578
rect 1119 16510 1237 16520
rect 1119 16448 1161 16510
rect 1195 16448 1237 16510
rect 1119 16442 1237 16448
rect 1119 16376 1161 16442
rect 1195 16376 1237 16442
rect 1119 16374 1237 16376
rect 1119 16340 1161 16374
rect 1195 16340 1237 16374
rect 1119 16338 1237 16340
rect 1119 16272 1161 16338
rect 1195 16272 1237 16338
rect 1119 16266 1237 16272
rect 1119 16204 1161 16266
rect 1195 16204 1237 16266
rect 1119 16194 1237 16204
rect 1119 16136 1161 16194
rect 1195 16136 1237 16194
rect 1119 16122 1237 16136
rect 1119 16068 1161 16122
rect 1195 16068 1237 16122
rect 1119 16050 1237 16068
rect 1119 16000 1161 16050
rect 1195 16000 1237 16050
rect 1119 15978 1237 16000
rect 1119 15932 1161 15978
rect 1195 15932 1237 15978
rect 1119 15906 1237 15932
rect 1119 15864 1161 15906
rect 1195 15864 1237 15906
rect 1119 15834 1237 15864
rect 1119 15796 1161 15834
rect 1195 15796 1237 15834
rect 1119 15762 1237 15796
rect 1119 15728 1161 15762
rect 1195 15728 1237 15762
rect 1119 15694 1237 15728
rect 1119 15656 1161 15694
rect 1195 15656 1237 15694
rect 1119 15626 1237 15656
rect 1119 15584 1161 15626
rect 1195 15584 1237 15626
rect 1119 15558 1237 15584
rect 1119 15512 1161 15558
rect 1195 15512 1237 15558
rect 1119 15490 1237 15512
rect 1119 15440 1161 15490
rect 1195 15440 1237 15490
rect 1119 15422 1237 15440
rect 1119 15368 1161 15422
rect 1195 15368 1237 15422
rect 1119 15319 1237 15368
rect 13769 24767 13809 24780
rect 13843 24767 13887 24801
rect 13769 24733 13887 24767
rect 13769 24699 13809 24733
rect 13843 24699 13887 24733
rect 13769 24665 13887 24699
rect 13769 24631 13809 24665
rect 13843 24631 13887 24665
rect 13769 24597 13887 24631
rect 13769 24563 13809 24597
rect 13843 24563 13887 24597
rect 13769 24529 13887 24563
rect 13769 24495 13809 24529
rect 13843 24495 13887 24529
rect 13769 24461 13887 24495
rect 13769 24427 13809 24461
rect 13843 24427 13887 24461
rect 13769 24393 13887 24427
rect 13769 24359 13809 24393
rect 13843 24359 13887 24393
rect 13769 24325 13887 24359
rect 13769 24291 13809 24325
rect 13843 24291 13887 24325
rect 13769 24257 13887 24291
rect 13769 24223 13809 24257
rect 13843 24223 13887 24257
rect 13769 24189 13887 24223
rect 13769 24155 13809 24189
rect 13843 24155 13887 24189
rect 13769 24121 13887 24155
rect 13769 24087 13809 24121
rect 13843 24087 13887 24121
rect 13769 24053 13887 24087
rect 13769 24019 13809 24053
rect 13843 24019 13887 24053
rect 13769 23985 13887 24019
rect 13769 23951 13809 23985
rect 13843 23951 13887 23985
rect 13769 23917 13887 23951
rect 13769 23883 13809 23917
rect 13843 23883 13887 23917
rect 13769 23849 13887 23883
rect 13769 23815 13809 23849
rect 13843 23815 13887 23849
rect 13769 23781 13887 23815
rect 13769 23747 13809 23781
rect 13843 23747 13887 23781
rect 13769 23713 13887 23747
rect 13769 23679 13809 23713
rect 13843 23679 13887 23713
rect 13769 23645 13887 23679
rect 13769 23611 13809 23645
rect 13843 23611 13887 23645
rect 13769 23577 13887 23611
rect 13769 23543 13809 23577
rect 13843 23543 13887 23577
rect 13769 23509 13887 23543
rect 13769 23475 13809 23509
rect 13843 23475 13887 23509
rect 13769 23441 13887 23475
rect 13769 23407 13809 23441
rect 13843 23407 13887 23441
rect 13769 23397 13887 23407
rect 13769 23339 13809 23397
rect 13843 23339 13887 23397
rect 13769 23325 13887 23339
rect 13769 23271 13809 23325
rect 13843 23271 13887 23325
rect 13769 23253 13887 23271
rect 13769 23203 13809 23253
rect 13843 23203 13887 23253
rect 13769 23181 13887 23203
rect 13769 23135 13809 23181
rect 13843 23135 13887 23181
rect 13769 23109 13887 23135
rect 13769 23067 13809 23109
rect 13843 23067 13887 23109
rect 13769 23037 13887 23067
rect 13769 22999 13809 23037
rect 13843 22999 13887 23037
rect 13769 22965 13887 22999
rect 13769 22931 13809 22965
rect 13843 22931 13887 22965
rect 13769 22897 13887 22931
rect 13769 22859 13809 22897
rect 13843 22859 13887 22897
rect 13769 22829 13887 22859
rect 13769 22787 13809 22829
rect 13843 22787 13887 22829
rect 13769 22761 13887 22787
rect 13769 22715 13809 22761
rect 13843 22715 13887 22761
rect 13769 22693 13887 22715
rect 13769 22643 13809 22693
rect 13843 22643 13887 22693
rect 13769 22625 13887 22643
rect 13769 22571 13809 22625
rect 13843 22571 13887 22625
rect 13769 22557 13887 22571
rect 13769 22499 13809 22557
rect 13843 22499 13887 22557
rect 13769 22489 13887 22499
rect 13769 22427 13809 22489
rect 13843 22427 13887 22489
rect 13769 22421 13887 22427
rect 13769 22355 13809 22421
rect 13843 22355 13887 22421
rect 13769 22353 13887 22355
rect 13769 22319 13809 22353
rect 13843 22319 13887 22353
rect 13769 22317 13887 22319
rect 13769 22251 13809 22317
rect 13843 22251 13887 22317
rect 13769 22245 13887 22251
rect 13769 22183 13809 22245
rect 13843 22183 13887 22245
rect 13769 22173 13887 22183
rect 13769 22115 13809 22173
rect 13843 22115 13887 22173
rect 13769 22101 13887 22115
rect 13769 22047 13809 22101
rect 13843 22047 13887 22101
rect 13769 22029 13887 22047
rect 13769 21979 13809 22029
rect 13843 21979 13887 22029
rect 13769 21957 13887 21979
rect 13769 21911 13809 21957
rect 13843 21911 13887 21957
rect 13769 21885 13887 21911
rect 13769 21843 13809 21885
rect 13843 21843 13887 21885
rect 13769 21813 13887 21843
rect 13769 21775 13809 21813
rect 13843 21775 13887 21813
rect 13769 21741 13887 21775
rect 13769 21707 13809 21741
rect 13843 21707 13887 21741
rect 13769 21673 13887 21707
rect 13769 21635 13809 21673
rect 13843 21635 13887 21673
rect 13769 21605 13887 21635
rect 13769 21563 13809 21605
rect 13843 21563 13887 21605
rect 13769 21537 13887 21563
rect 13769 21491 13809 21537
rect 13843 21491 13887 21537
rect 13769 21469 13887 21491
rect 13769 21419 13809 21469
rect 13843 21419 13887 21469
rect 13769 21401 13887 21419
rect 13769 21347 13809 21401
rect 13843 21347 13887 21401
rect 13769 21333 13887 21347
rect 13769 21275 13809 21333
rect 13843 21275 13887 21333
rect 13769 21265 13887 21275
rect 13769 21203 13809 21265
rect 13843 21203 13887 21265
rect 13769 21197 13887 21203
rect 13769 21131 13809 21197
rect 13843 21131 13887 21197
rect 13769 21129 13887 21131
rect 13769 21095 13809 21129
rect 13843 21095 13887 21129
rect 13769 21093 13887 21095
rect 13769 21027 13809 21093
rect 13843 21027 13887 21093
rect 13769 21021 13887 21027
rect 13769 20959 13809 21021
rect 13843 20959 13887 21021
rect 13769 20949 13887 20959
rect 13769 20891 13809 20949
rect 13843 20891 13887 20949
rect 13769 20877 13887 20891
rect 13769 20823 13809 20877
rect 13843 20823 13887 20877
rect 13769 20805 13887 20823
rect 13769 20755 13809 20805
rect 13843 20755 13887 20805
rect 13769 20733 13887 20755
rect 13769 20687 13809 20733
rect 13843 20687 13887 20733
rect 13769 20661 13887 20687
rect 13769 20619 13809 20661
rect 13843 20619 13887 20661
rect 13769 20589 13887 20619
rect 13769 20551 13809 20589
rect 13843 20551 13887 20589
rect 13769 20517 13887 20551
rect 13769 20483 13809 20517
rect 13843 20483 13887 20517
rect 13769 20449 13887 20483
rect 13769 20411 13809 20449
rect 13843 20411 13887 20449
rect 13769 20381 13887 20411
rect 13769 20339 13809 20381
rect 13843 20339 13887 20381
rect 13769 20313 13887 20339
rect 13769 20267 13809 20313
rect 13843 20267 13887 20313
rect 13769 20245 13887 20267
rect 13769 20195 13809 20245
rect 13843 20195 13887 20245
rect 13769 20177 13887 20195
rect 13769 20123 13809 20177
rect 13843 20123 13887 20177
rect 13769 20109 13887 20123
rect 13769 20051 13809 20109
rect 13843 20051 13887 20109
rect 13769 20041 13887 20051
rect 13769 19979 13809 20041
rect 13843 19979 13887 20041
rect 13769 19973 13887 19979
rect 13769 19907 13809 19973
rect 13843 19907 13887 19973
rect 13769 19905 13887 19907
rect 13769 19871 13809 19905
rect 13843 19871 13887 19905
rect 13769 19869 13887 19871
rect 13769 19803 13809 19869
rect 13843 19803 13887 19869
rect 13769 19797 13887 19803
rect 13769 19735 13809 19797
rect 13843 19735 13887 19797
rect 13769 19725 13887 19735
rect 13769 19667 13809 19725
rect 13843 19667 13887 19725
rect 13769 19653 13887 19667
rect 13769 19599 13809 19653
rect 13843 19599 13887 19653
rect 13769 19581 13887 19599
rect 13769 19531 13809 19581
rect 13843 19531 13887 19581
rect 13769 19509 13887 19531
rect 13769 19463 13809 19509
rect 13843 19463 13887 19509
rect 13769 19437 13887 19463
rect 13769 19395 13809 19437
rect 13843 19395 13887 19437
rect 13769 19365 13887 19395
rect 13769 19327 13809 19365
rect 13843 19327 13887 19365
rect 13769 19293 13887 19327
rect 13769 19259 13809 19293
rect 13843 19259 13887 19293
rect 13769 19225 13887 19259
rect 13769 19187 13809 19225
rect 13843 19187 13887 19225
rect 13769 19157 13887 19187
rect 13769 19115 13809 19157
rect 13843 19115 13887 19157
rect 13769 19089 13887 19115
rect 13769 19043 13809 19089
rect 13843 19043 13887 19089
rect 13769 19021 13887 19043
rect 13769 18971 13809 19021
rect 13843 18971 13887 19021
rect 13769 18953 13887 18971
rect 13769 18899 13809 18953
rect 13843 18899 13887 18953
rect 13769 18885 13887 18899
rect 13769 18827 13809 18885
rect 13843 18827 13887 18885
rect 13769 18817 13887 18827
rect 13769 18755 13809 18817
rect 13843 18755 13887 18817
rect 13769 18749 13887 18755
rect 13769 18683 13809 18749
rect 13843 18683 13887 18749
rect 13769 18681 13887 18683
rect 13769 18647 13809 18681
rect 13843 18647 13887 18681
rect 13769 18645 13887 18647
rect 13769 18579 13809 18645
rect 13843 18579 13887 18645
rect 13769 18573 13887 18579
rect 13769 18511 13809 18573
rect 13843 18511 13887 18573
rect 13769 18501 13887 18511
rect 13769 18443 13809 18501
rect 13843 18443 13887 18501
rect 13769 18429 13887 18443
rect 13769 18375 13809 18429
rect 13843 18375 13887 18429
rect 13769 18357 13887 18375
rect 13769 18307 13809 18357
rect 13843 18307 13887 18357
rect 13769 18285 13887 18307
rect 13769 18239 13809 18285
rect 13843 18239 13887 18285
rect 13769 18213 13887 18239
rect 13769 18171 13809 18213
rect 13843 18171 13887 18213
rect 13769 18141 13887 18171
rect 13769 18103 13809 18141
rect 13843 18103 13887 18141
rect 13769 18069 13887 18103
rect 13769 18035 13809 18069
rect 13843 18035 13887 18069
rect 13769 18001 13887 18035
rect 13769 17963 13809 18001
rect 13843 17963 13887 18001
rect 13769 17933 13887 17963
rect 13769 17891 13809 17933
rect 13843 17891 13887 17933
rect 13769 17865 13887 17891
rect 13769 17819 13809 17865
rect 13843 17819 13887 17865
rect 13769 17797 13887 17819
rect 13769 17747 13809 17797
rect 13843 17747 13887 17797
rect 13769 17729 13887 17747
rect 13769 17675 13809 17729
rect 13843 17675 13887 17729
rect 13769 17661 13887 17675
rect 13769 17603 13809 17661
rect 13843 17603 13887 17661
rect 13769 17593 13887 17603
rect 13769 17531 13809 17593
rect 13843 17531 13887 17593
rect 13769 17525 13887 17531
rect 13769 17459 13809 17525
rect 13843 17459 13887 17525
rect 13769 17457 13887 17459
rect 13769 17423 13809 17457
rect 13843 17423 13887 17457
rect 13769 17421 13887 17423
rect 13769 17355 13809 17421
rect 13843 17355 13887 17421
rect 13769 17349 13887 17355
rect 13769 17287 13809 17349
rect 13843 17287 13887 17349
rect 13769 17277 13887 17287
rect 13769 17219 13809 17277
rect 13843 17219 13887 17277
rect 13769 17205 13887 17219
rect 13769 17151 13809 17205
rect 13843 17151 13887 17205
rect 13769 17133 13887 17151
rect 13769 17083 13809 17133
rect 13843 17083 13887 17133
rect 13769 17061 13887 17083
rect 13769 17015 13809 17061
rect 13843 17015 13887 17061
rect 13769 16989 13887 17015
rect 13769 16947 13809 16989
rect 13843 16947 13887 16989
rect 13769 16917 13887 16947
rect 13769 16879 13809 16917
rect 13843 16879 13887 16917
rect 13769 16845 13887 16879
rect 13769 16811 13809 16845
rect 13843 16811 13887 16845
rect 13769 16777 13887 16811
rect 13769 16739 13809 16777
rect 13843 16739 13887 16777
rect 13769 16709 13887 16739
rect 13769 16667 13809 16709
rect 13843 16667 13887 16709
rect 13769 16641 13887 16667
rect 13769 16595 13809 16641
rect 13843 16595 13887 16641
rect 13769 16573 13887 16595
rect 13769 16523 13809 16573
rect 13843 16523 13887 16573
rect 13769 16505 13887 16523
rect 13769 16451 13809 16505
rect 13843 16451 13887 16505
rect 13769 16437 13887 16451
rect 13769 16379 13809 16437
rect 13843 16379 13887 16437
rect 13769 16369 13887 16379
rect 13769 16307 13809 16369
rect 13843 16307 13887 16369
rect 13769 16301 13887 16307
rect 13769 16235 13809 16301
rect 13843 16235 13887 16301
rect 13769 16233 13887 16235
rect 13769 16199 13809 16233
rect 13843 16199 13887 16233
rect 13769 16197 13887 16199
rect 13769 16131 13809 16197
rect 13843 16131 13887 16197
rect 13769 16125 13887 16131
rect 13769 16063 13809 16125
rect 13843 16063 13887 16125
rect 13769 16053 13887 16063
rect 13769 15995 13809 16053
rect 13843 15995 13887 16053
rect 13769 15981 13887 15995
rect 13769 15927 13809 15981
rect 13843 15927 13887 15981
rect 13769 15909 13887 15927
rect 13769 15859 13809 15909
rect 13843 15859 13887 15909
rect 13769 15837 13887 15859
rect 13769 15791 13809 15837
rect 13843 15791 13887 15837
rect 13769 15765 13887 15791
rect 13769 15723 13809 15765
rect 13843 15723 13887 15765
rect 13769 15693 13887 15723
rect 13769 15655 13809 15693
rect 13843 15655 13887 15693
rect 13769 15621 13887 15655
rect 13769 15587 13809 15621
rect 13843 15587 13887 15621
rect 13769 15553 13887 15587
rect 13769 15515 13809 15553
rect 13843 15515 13887 15553
rect 13769 15485 13887 15515
rect 13769 15443 13809 15485
rect 13843 15443 13887 15485
rect 13769 15417 13887 15443
rect 13769 15371 13809 15417
rect 13843 15371 13887 15417
rect 13769 15319 13887 15371
rect 1119 15278 13887 15319
rect 1119 15244 1298 15278
rect 1336 15244 1370 15278
rect 1404 15244 1438 15278
rect 1476 15244 1506 15278
rect 1548 15244 1574 15278
rect 1620 15244 1642 15278
rect 1692 15244 1710 15278
rect 1764 15244 1778 15278
rect 1836 15244 1846 15278
rect 1908 15244 1914 15278
rect 1980 15244 1982 15278
rect 2016 15244 2018 15278
rect 2084 15244 2090 15278
rect 2152 15244 2162 15278
rect 2220 15244 2234 15278
rect 2288 15244 2306 15278
rect 2356 15244 2378 15278
rect 2424 15244 2450 15278
rect 2492 15244 2522 15278
rect 2560 15244 2594 15278
rect 2628 15244 2662 15278
rect 2700 15244 2730 15278
rect 2772 15244 2798 15278
rect 2844 15244 2866 15278
rect 2916 15244 2934 15278
rect 2988 15244 3002 15278
rect 3060 15244 3070 15278
rect 3132 15244 3138 15278
rect 3204 15244 3206 15278
rect 3240 15244 3242 15278
rect 3308 15244 3314 15278
rect 3376 15244 3386 15278
rect 3444 15244 3458 15278
rect 3512 15244 3530 15278
rect 3580 15244 3602 15278
rect 3648 15244 3674 15278
rect 3716 15244 3746 15278
rect 3784 15244 3818 15278
rect 3852 15244 3886 15278
rect 3924 15244 3954 15278
rect 3996 15244 4022 15278
rect 4068 15244 4090 15278
rect 4140 15244 4158 15278
rect 4212 15244 4226 15278
rect 4284 15244 4294 15278
rect 4356 15244 4362 15278
rect 4428 15244 4430 15278
rect 4464 15244 4466 15278
rect 4532 15244 4538 15278
rect 4600 15244 4610 15278
rect 4668 15244 4682 15278
rect 4736 15244 4754 15278
rect 4804 15244 4826 15278
rect 4872 15244 4898 15278
rect 4940 15244 4970 15278
rect 5008 15244 5042 15278
rect 5076 15244 5110 15278
rect 5148 15244 5178 15278
rect 5220 15244 5246 15278
rect 5292 15244 5314 15278
rect 5364 15244 5382 15278
rect 5436 15244 5450 15278
rect 5508 15244 5518 15278
rect 5580 15244 5586 15278
rect 5652 15244 5654 15278
rect 5688 15244 5690 15278
rect 5756 15244 5762 15278
rect 5824 15244 5834 15278
rect 5892 15244 5906 15278
rect 5960 15244 5978 15278
rect 6028 15244 6050 15278
rect 6096 15244 6122 15278
rect 6164 15244 6194 15278
rect 6232 15244 6266 15278
rect 6300 15244 6334 15278
rect 6372 15244 6402 15278
rect 6444 15244 6470 15278
rect 6516 15244 6538 15278
rect 6588 15244 6606 15278
rect 6660 15244 6674 15278
rect 6732 15244 6742 15278
rect 6804 15244 6810 15278
rect 6876 15244 6878 15278
rect 6912 15244 6914 15278
rect 6980 15244 6986 15278
rect 7048 15244 7058 15278
rect 7116 15244 7130 15278
rect 7184 15244 7202 15278
rect 7252 15244 7274 15278
rect 7320 15244 7346 15278
rect 7388 15244 7418 15278
rect 7456 15244 7490 15278
rect 7524 15244 7558 15278
rect 7596 15244 7626 15278
rect 7668 15244 7694 15278
rect 7740 15244 7762 15278
rect 7812 15244 7830 15278
rect 7884 15244 7898 15278
rect 7956 15244 7966 15278
rect 8028 15244 8034 15278
rect 8100 15244 8102 15278
rect 8136 15244 8138 15278
rect 8204 15244 8210 15278
rect 8272 15244 8282 15278
rect 8340 15244 8354 15278
rect 8408 15244 8426 15278
rect 8476 15244 8498 15278
rect 8544 15244 8570 15278
rect 8612 15244 8642 15278
rect 8680 15244 8714 15278
rect 8748 15244 8782 15278
rect 8820 15244 8850 15278
rect 8892 15244 8918 15278
rect 8964 15244 8986 15278
rect 9036 15244 9054 15278
rect 9108 15244 9122 15278
rect 9180 15244 9190 15278
rect 9252 15244 9258 15278
rect 9324 15244 9326 15278
rect 9360 15244 9362 15278
rect 9428 15244 9434 15278
rect 9496 15244 9506 15278
rect 9564 15244 9578 15278
rect 9632 15244 9650 15278
rect 9700 15244 9722 15278
rect 9768 15244 9794 15278
rect 9836 15244 9866 15278
rect 9904 15244 9938 15278
rect 9972 15244 10006 15278
rect 10044 15244 10074 15278
rect 10116 15244 10142 15278
rect 10188 15244 10210 15278
rect 10260 15244 10278 15278
rect 10332 15244 10346 15278
rect 10404 15244 10414 15278
rect 10476 15244 10482 15278
rect 10548 15244 10550 15278
rect 10584 15244 10586 15278
rect 10652 15244 10658 15278
rect 10720 15244 10730 15278
rect 10788 15244 10802 15278
rect 10856 15244 10874 15278
rect 10924 15244 10946 15278
rect 10992 15244 11018 15278
rect 11060 15244 11090 15278
rect 11128 15244 11162 15278
rect 11196 15244 11230 15278
rect 11268 15244 11298 15278
rect 11340 15244 11366 15278
rect 11412 15244 11434 15278
rect 11484 15244 11502 15278
rect 11556 15244 11570 15278
rect 11628 15244 11638 15278
rect 11700 15244 11706 15278
rect 11772 15244 11774 15278
rect 11808 15244 11810 15278
rect 11876 15244 11882 15278
rect 11944 15244 11954 15278
rect 12012 15244 12026 15278
rect 12080 15244 12098 15278
rect 12148 15244 12170 15278
rect 12216 15244 12242 15278
rect 12284 15244 12314 15278
rect 12352 15244 12386 15278
rect 12420 15244 12454 15278
rect 12492 15244 12522 15278
rect 12564 15244 12590 15278
rect 12636 15244 12658 15278
rect 12708 15244 12726 15278
rect 12780 15244 12794 15278
rect 12852 15244 12862 15278
rect 12924 15244 12930 15278
rect 12996 15244 12998 15278
rect 13032 15244 13034 15278
rect 13100 15244 13106 15278
rect 13168 15244 13178 15278
rect 13236 15244 13250 15278
rect 13304 15244 13322 15278
rect 13372 15244 13394 15278
rect 13440 15244 13466 15278
rect 13508 15244 13538 15278
rect 13576 15244 13610 15278
rect 13644 15244 13678 15278
rect 13716 15244 13887 15278
rect 1119 15201 13887 15244
rect 13968 34707 14122 34741
rect 14156 34724 14297 34741
rect 14331 34724 14361 34758
rect 14156 34707 14361 34724
rect 13968 34690 14361 34707
rect 13968 34669 14297 34690
rect 13968 34635 14122 34669
rect 14156 34656 14297 34669
rect 14331 34656 14361 34690
rect 14156 34635 14361 34656
rect 13968 34622 14361 34635
rect 13968 34597 14297 34622
rect 13968 34563 14122 34597
rect 14156 34588 14297 34597
rect 14331 34588 14361 34622
rect 14156 34563 14361 34588
rect 13968 34554 14361 34563
rect 13968 34525 14297 34554
rect 13968 34491 14122 34525
rect 14156 34520 14297 34525
rect 14331 34520 14361 34554
rect 14156 34491 14361 34520
rect 13968 34486 14361 34491
rect 13968 34453 14297 34486
rect 13968 34419 14122 34453
rect 14156 34452 14297 34453
rect 14331 34452 14361 34486
rect 14156 34419 14361 34452
rect 13968 34418 14361 34419
rect 13968 34384 14297 34418
rect 14331 34384 14361 34418
rect 13968 34381 14361 34384
rect 13968 34347 14122 34381
rect 14156 34350 14361 34381
rect 14156 34347 14297 34350
rect 13968 34316 14297 34347
rect 14331 34316 14361 34350
rect 13968 34309 14361 34316
rect 13968 34275 14122 34309
rect 14156 34282 14361 34309
rect 14156 34275 14297 34282
rect 13968 34248 14297 34275
rect 14331 34248 14361 34282
rect 13968 34237 14361 34248
rect 13968 34203 14122 34237
rect 14156 34214 14361 34237
rect 14156 34203 14297 34214
rect 13968 34180 14297 34203
rect 14331 34180 14361 34214
rect 13968 34165 14361 34180
rect 13968 34131 14122 34165
rect 14156 34146 14361 34165
rect 14156 34131 14297 34146
rect 13968 34112 14297 34131
rect 14331 34112 14361 34146
rect 13968 34093 14361 34112
rect 13968 34059 14122 34093
rect 14156 34078 14361 34093
rect 14156 34059 14297 34078
rect 13968 34044 14297 34059
rect 14331 34044 14361 34078
rect 13968 34021 14361 34044
rect 13968 33987 14122 34021
rect 14156 34010 14361 34021
rect 14156 33987 14297 34010
rect 13968 33976 14297 33987
rect 14331 33976 14361 34010
rect 13968 33949 14361 33976
rect 13968 33915 14122 33949
rect 14156 33942 14361 33949
rect 14156 33915 14297 33942
rect 13968 33908 14297 33915
rect 14331 33908 14361 33942
rect 13968 33877 14361 33908
rect 13968 33843 14122 33877
rect 14156 33874 14361 33877
rect 14156 33843 14297 33874
rect 13968 33840 14297 33843
rect 14331 33840 14361 33874
rect 13968 33806 14361 33840
rect 13968 33805 14297 33806
rect 13968 33771 14122 33805
rect 14156 33772 14297 33805
rect 14331 33772 14361 33806
rect 14156 33771 14361 33772
rect 13968 33738 14361 33771
rect 13968 33733 14297 33738
rect 13968 33699 14122 33733
rect 14156 33704 14297 33733
rect 14331 33704 14361 33738
rect 14156 33699 14361 33704
rect 13968 33670 14361 33699
rect 13968 33661 14297 33670
rect 13968 33627 14122 33661
rect 14156 33636 14297 33661
rect 14331 33636 14361 33670
rect 14156 33627 14361 33636
rect 13968 33602 14361 33627
rect 13968 33589 14297 33602
rect 13968 33555 14122 33589
rect 14156 33568 14297 33589
rect 14331 33568 14361 33602
rect 14156 33555 14361 33568
rect 13968 33534 14361 33555
rect 13968 33517 14297 33534
rect 13968 33483 14122 33517
rect 14156 33500 14297 33517
rect 14331 33500 14361 33534
rect 14156 33483 14361 33500
rect 13968 33466 14361 33483
rect 13968 33445 14297 33466
rect 13968 33411 14122 33445
rect 14156 33432 14297 33445
rect 14331 33432 14361 33466
rect 14156 33411 14361 33432
rect 13968 33398 14361 33411
rect 13968 33373 14297 33398
rect 13968 33339 14122 33373
rect 14156 33364 14297 33373
rect 14331 33364 14361 33398
rect 14156 33339 14361 33364
rect 13968 33330 14361 33339
rect 13968 33301 14297 33330
rect 13968 33267 14122 33301
rect 14156 33296 14297 33301
rect 14331 33296 14361 33330
rect 14156 33267 14361 33296
rect 13968 33262 14361 33267
rect 13968 33229 14297 33262
rect 13968 33195 14122 33229
rect 14156 33228 14297 33229
rect 14331 33228 14361 33262
rect 14156 33195 14361 33228
rect 13968 33194 14361 33195
rect 13968 33160 14297 33194
rect 14331 33160 14361 33194
rect 13968 33157 14361 33160
rect 13968 33123 14122 33157
rect 14156 33126 14361 33157
rect 14156 33123 14297 33126
rect 13968 33092 14297 33123
rect 14331 33092 14361 33126
rect 13968 33085 14361 33092
rect 13968 33051 14122 33085
rect 14156 33058 14361 33085
rect 14156 33051 14297 33058
rect 13968 33024 14297 33051
rect 14331 33024 14361 33058
rect 13968 33013 14361 33024
rect 13968 32979 14122 33013
rect 14156 32990 14361 33013
rect 14156 32979 14297 32990
rect 13968 32956 14297 32979
rect 14331 32956 14361 32990
rect 13968 32941 14361 32956
rect 13968 32907 14122 32941
rect 14156 32922 14361 32941
rect 14156 32907 14297 32922
rect 13968 32888 14297 32907
rect 14331 32888 14361 32922
rect 13968 32869 14361 32888
rect 13968 32835 14122 32869
rect 14156 32854 14361 32869
rect 14156 32835 14297 32854
rect 13968 32820 14297 32835
rect 14331 32820 14361 32854
rect 13968 32797 14361 32820
rect 13968 32763 14122 32797
rect 14156 32786 14361 32797
rect 14156 32763 14297 32786
rect 13968 32752 14297 32763
rect 14331 32752 14361 32786
rect 13968 32725 14361 32752
rect 13968 32691 14122 32725
rect 14156 32718 14361 32725
rect 14156 32691 14297 32718
rect 13968 32684 14297 32691
rect 14331 32684 14361 32718
rect 13968 32653 14361 32684
rect 13968 32619 14122 32653
rect 14156 32650 14361 32653
rect 14156 32619 14297 32650
rect 13968 32616 14297 32619
rect 14331 32616 14361 32650
rect 13968 32582 14361 32616
rect 13968 32581 14297 32582
rect 13968 32547 14122 32581
rect 14156 32548 14297 32581
rect 14331 32548 14361 32582
rect 14156 32547 14361 32548
rect 13968 32514 14361 32547
rect 13968 32509 14297 32514
rect 13968 32475 14122 32509
rect 14156 32480 14297 32509
rect 14331 32480 14361 32514
rect 14156 32475 14361 32480
rect 13968 32446 14361 32475
rect 13968 32437 14297 32446
rect 13968 32403 14122 32437
rect 14156 32412 14297 32437
rect 14331 32412 14361 32446
rect 14156 32403 14361 32412
rect 13968 32378 14361 32403
rect 13968 32365 14297 32378
rect 13968 32331 14122 32365
rect 14156 32344 14297 32365
rect 14331 32344 14361 32378
rect 14156 32331 14361 32344
rect 13968 32310 14361 32331
rect 13968 32293 14297 32310
rect 13968 32259 14122 32293
rect 14156 32276 14297 32293
rect 14331 32276 14361 32310
rect 14156 32259 14361 32276
rect 13968 32242 14361 32259
rect 13968 32221 14297 32242
rect 13968 32187 14122 32221
rect 14156 32208 14297 32221
rect 14331 32208 14361 32242
rect 14156 32187 14361 32208
rect 13968 32174 14361 32187
rect 13968 32149 14297 32174
rect 13968 32115 14122 32149
rect 14156 32140 14297 32149
rect 14331 32140 14361 32174
rect 14156 32115 14361 32140
rect 13968 32106 14361 32115
rect 13968 32077 14297 32106
rect 13968 32043 14122 32077
rect 14156 32072 14297 32077
rect 14331 32072 14361 32106
rect 14156 32043 14361 32072
rect 13968 32038 14361 32043
rect 13968 32005 14297 32038
rect 13968 31971 14122 32005
rect 14156 32004 14297 32005
rect 14331 32004 14361 32038
rect 14156 31971 14361 32004
rect 13968 31970 14361 31971
rect 13968 31936 14297 31970
rect 14331 31936 14361 31970
rect 13968 31933 14361 31936
rect 13968 31899 14122 31933
rect 14156 31902 14361 31933
rect 14156 31899 14297 31902
rect 13968 31868 14297 31899
rect 14331 31868 14361 31902
rect 13968 31861 14361 31868
rect 13968 31827 14122 31861
rect 14156 31834 14361 31861
rect 14156 31827 14297 31834
rect 13968 31800 14297 31827
rect 14331 31800 14361 31834
rect 13968 31789 14361 31800
rect 13968 31755 14122 31789
rect 14156 31766 14361 31789
rect 14156 31755 14297 31766
rect 13968 31732 14297 31755
rect 14331 31732 14361 31766
rect 13968 31717 14361 31732
rect 13968 31683 14122 31717
rect 14156 31698 14361 31717
rect 14156 31683 14297 31698
rect 13968 31664 14297 31683
rect 14331 31664 14361 31698
rect 13968 31645 14361 31664
rect 13968 31611 14122 31645
rect 14156 31630 14361 31645
rect 14156 31611 14297 31630
rect 13968 31596 14297 31611
rect 14331 31596 14361 31630
rect 13968 31573 14361 31596
rect 13968 31539 14122 31573
rect 14156 31562 14361 31573
rect 14156 31539 14297 31562
rect 13968 31528 14297 31539
rect 14331 31528 14361 31562
rect 13968 31501 14361 31528
rect 13968 31467 14122 31501
rect 14156 31494 14361 31501
rect 14156 31467 14297 31494
rect 13968 31460 14297 31467
rect 14331 31460 14361 31494
rect 13968 31429 14361 31460
rect 13968 31395 14122 31429
rect 14156 31426 14361 31429
rect 14156 31395 14297 31426
rect 13968 31392 14297 31395
rect 14331 31392 14361 31426
rect 13968 31358 14361 31392
rect 13968 31357 14297 31358
rect 13968 31323 14122 31357
rect 14156 31324 14297 31357
rect 14331 31324 14361 31358
rect 14156 31323 14361 31324
rect 13968 31290 14361 31323
rect 13968 31285 14297 31290
rect 13968 31251 14122 31285
rect 14156 31256 14297 31285
rect 14331 31256 14361 31290
rect 14156 31251 14361 31256
rect 13968 31222 14361 31251
rect 13968 31213 14297 31222
rect 13968 31179 14122 31213
rect 14156 31188 14297 31213
rect 14331 31188 14361 31222
rect 14156 31179 14361 31188
rect 13968 31154 14361 31179
rect 13968 31141 14297 31154
rect 13968 31107 14122 31141
rect 14156 31120 14297 31141
rect 14331 31120 14361 31154
rect 14156 31107 14361 31120
rect 13968 31086 14361 31107
rect 13968 31069 14297 31086
rect 13968 31035 14122 31069
rect 14156 31052 14297 31069
rect 14331 31052 14361 31086
rect 14156 31035 14361 31052
rect 13968 31018 14361 31035
rect 13968 30997 14297 31018
rect 13968 30963 14122 30997
rect 14156 30984 14297 30997
rect 14331 30984 14361 31018
rect 14156 30963 14361 30984
rect 13968 30950 14361 30963
rect 13968 30925 14297 30950
rect 13968 30891 14122 30925
rect 14156 30916 14297 30925
rect 14331 30916 14361 30950
rect 14156 30891 14361 30916
rect 13968 30882 14361 30891
rect 13968 30853 14297 30882
rect 13968 30819 14122 30853
rect 14156 30848 14297 30853
rect 14331 30848 14361 30882
rect 14156 30819 14361 30848
rect 13968 30814 14361 30819
rect 13968 30781 14297 30814
rect 13968 30747 14122 30781
rect 14156 30780 14297 30781
rect 14331 30780 14361 30814
rect 14156 30747 14361 30780
rect 13968 30746 14361 30747
rect 13968 30712 14297 30746
rect 14331 30712 14361 30746
rect 13968 30709 14361 30712
rect 13968 30675 14122 30709
rect 14156 30678 14361 30709
rect 14156 30675 14297 30678
rect 13968 30644 14297 30675
rect 14331 30644 14361 30678
rect 13968 30637 14361 30644
rect 13968 30603 14122 30637
rect 14156 30610 14361 30637
rect 14156 30603 14297 30610
rect 13968 30576 14297 30603
rect 14331 30576 14361 30610
rect 13968 30565 14361 30576
rect 13968 30531 14122 30565
rect 14156 30542 14361 30565
rect 14156 30531 14297 30542
rect 13968 30508 14297 30531
rect 14331 30508 14361 30542
rect 13968 30493 14361 30508
rect 13968 30459 14122 30493
rect 14156 30474 14361 30493
rect 14156 30459 14297 30474
rect 13968 30440 14297 30459
rect 14331 30440 14361 30474
rect 13968 30421 14361 30440
rect 13968 30387 14122 30421
rect 14156 30406 14361 30421
rect 14156 30387 14297 30406
rect 13968 30372 14297 30387
rect 14331 30372 14361 30406
rect 13968 30349 14361 30372
rect 13968 30315 14122 30349
rect 14156 30338 14361 30349
rect 14156 30315 14297 30338
rect 13968 30304 14297 30315
rect 14331 30304 14361 30338
rect 13968 30277 14361 30304
rect 13968 30243 14122 30277
rect 14156 30270 14361 30277
rect 14156 30243 14297 30270
rect 13968 30236 14297 30243
rect 14331 30236 14361 30270
rect 13968 30205 14361 30236
rect 13968 30171 14122 30205
rect 14156 30202 14361 30205
rect 14156 30171 14297 30202
rect 13968 30168 14297 30171
rect 14331 30168 14361 30202
rect 13968 30134 14361 30168
rect 13968 30133 14297 30134
rect 13968 30099 14122 30133
rect 14156 30100 14297 30133
rect 14331 30100 14361 30134
rect 14156 30099 14361 30100
rect 13968 30066 14361 30099
rect 13968 30061 14297 30066
rect 13968 30027 14122 30061
rect 14156 30032 14297 30061
rect 14331 30032 14361 30066
rect 14156 30027 14361 30032
rect 13968 29998 14361 30027
rect 13968 29989 14297 29998
rect 13968 29955 14122 29989
rect 14156 29964 14297 29989
rect 14331 29964 14361 29998
rect 14156 29955 14361 29964
rect 13968 29930 14361 29955
rect 13968 29917 14297 29930
rect 13968 29883 14122 29917
rect 14156 29896 14297 29917
rect 14331 29896 14361 29930
rect 14156 29883 14361 29896
rect 13968 29862 14361 29883
rect 13968 29845 14297 29862
rect 13968 29811 14122 29845
rect 14156 29828 14297 29845
rect 14331 29828 14361 29862
rect 14156 29811 14361 29828
rect 13968 29794 14361 29811
rect 13968 29773 14297 29794
rect 13968 29739 14122 29773
rect 14156 29760 14297 29773
rect 14331 29760 14361 29794
rect 14156 29739 14361 29760
rect 13968 29726 14361 29739
rect 13968 29701 14297 29726
rect 13968 29667 14122 29701
rect 14156 29692 14297 29701
rect 14331 29692 14361 29726
rect 14156 29667 14361 29692
rect 13968 29658 14361 29667
rect 13968 29629 14297 29658
rect 13968 29595 14122 29629
rect 14156 29624 14297 29629
rect 14331 29624 14361 29658
rect 14156 29595 14361 29624
rect 13968 29590 14361 29595
rect 13968 29557 14297 29590
rect 13968 29523 14122 29557
rect 14156 29556 14297 29557
rect 14331 29556 14361 29590
rect 14156 29523 14361 29556
rect 13968 29522 14361 29523
rect 13968 29488 14297 29522
rect 14331 29488 14361 29522
rect 13968 29485 14361 29488
rect 13968 29451 14122 29485
rect 14156 29454 14361 29485
rect 14156 29451 14297 29454
rect 13968 29420 14297 29451
rect 14331 29420 14361 29454
rect 13968 29413 14361 29420
rect 13968 29379 14122 29413
rect 14156 29386 14361 29413
rect 14156 29379 14297 29386
rect 13968 29352 14297 29379
rect 14331 29352 14361 29386
rect 13968 29341 14361 29352
rect 13968 29307 14122 29341
rect 14156 29318 14361 29341
rect 14156 29307 14297 29318
rect 13968 29284 14297 29307
rect 14331 29284 14361 29318
rect 13968 29269 14361 29284
rect 13968 29235 14122 29269
rect 14156 29250 14361 29269
rect 14156 29235 14297 29250
rect 13968 29216 14297 29235
rect 14331 29216 14361 29250
rect 13968 29197 14361 29216
rect 13968 29163 14122 29197
rect 14156 29182 14361 29197
rect 14156 29163 14297 29182
rect 13968 29148 14297 29163
rect 14331 29148 14361 29182
rect 13968 29125 14361 29148
rect 13968 29091 14122 29125
rect 14156 29114 14361 29125
rect 14156 29091 14297 29114
rect 13968 29080 14297 29091
rect 14331 29080 14361 29114
rect 13968 29053 14361 29080
rect 13968 29019 14122 29053
rect 14156 29046 14361 29053
rect 14156 29019 14297 29046
rect 13968 29012 14297 29019
rect 14331 29012 14361 29046
rect 13968 28981 14361 29012
rect 13968 28947 14122 28981
rect 14156 28978 14361 28981
rect 14156 28947 14297 28978
rect 13968 28944 14297 28947
rect 14331 28944 14361 28978
rect 13968 28910 14361 28944
rect 13968 28909 14297 28910
rect 13968 28875 14122 28909
rect 14156 28876 14297 28909
rect 14331 28876 14361 28910
rect 14156 28875 14361 28876
rect 13968 28842 14361 28875
rect 13968 28837 14297 28842
rect 13968 28803 14122 28837
rect 14156 28808 14297 28837
rect 14331 28808 14361 28842
rect 14156 28803 14361 28808
rect 13968 28774 14361 28803
rect 13968 28765 14297 28774
rect 13968 28731 14122 28765
rect 14156 28740 14297 28765
rect 14331 28740 14361 28774
rect 14156 28731 14361 28740
rect 13968 28706 14361 28731
rect 13968 28693 14297 28706
rect 13968 28659 14122 28693
rect 14156 28672 14297 28693
rect 14331 28672 14361 28706
rect 14156 28659 14361 28672
rect 13968 28638 14361 28659
rect 13968 28621 14297 28638
rect 13968 28587 14122 28621
rect 14156 28604 14297 28621
rect 14331 28604 14361 28638
rect 14156 28587 14361 28604
rect 13968 28570 14361 28587
rect 13968 28549 14297 28570
rect 13968 28515 14122 28549
rect 14156 28536 14297 28549
rect 14331 28536 14361 28570
rect 14156 28515 14361 28536
rect 13968 28502 14361 28515
rect 13968 28477 14297 28502
rect 13968 28443 14122 28477
rect 14156 28468 14297 28477
rect 14331 28468 14361 28502
rect 14156 28443 14361 28468
rect 13968 28434 14361 28443
rect 13968 28405 14297 28434
rect 13968 28371 14122 28405
rect 14156 28400 14297 28405
rect 14331 28400 14361 28434
rect 14156 28371 14361 28400
rect 13968 28366 14361 28371
rect 13968 28333 14297 28366
rect 13968 28299 14122 28333
rect 14156 28332 14297 28333
rect 14331 28332 14361 28366
rect 14156 28299 14361 28332
rect 13968 28298 14361 28299
rect 13968 28264 14297 28298
rect 14331 28264 14361 28298
rect 13968 28261 14361 28264
rect 13968 28227 14122 28261
rect 14156 28230 14361 28261
rect 14156 28227 14297 28230
rect 13968 28196 14297 28227
rect 14331 28196 14361 28230
rect 13968 28189 14361 28196
rect 13968 28155 14122 28189
rect 14156 28162 14361 28189
rect 14156 28155 14297 28162
rect 13968 28128 14297 28155
rect 14331 28128 14361 28162
rect 13968 28117 14361 28128
rect 13968 28083 14122 28117
rect 14156 28094 14361 28117
rect 14156 28083 14297 28094
rect 13968 28060 14297 28083
rect 14331 28060 14361 28094
rect 13968 28045 14361 28060
rect 13968 28011 14122 28045
rect 14156 28026 14361 28045
rect 14156 28011 14297 28026
rect 13968 27992 14297 28011
rect 14331 27992 14361 28026
rect 13968 27973 14361 27992
rect 13968 27939 14122 27973
rect 14156 27958 14361 27973
rect 14156 27939 14297 27958
rect 13968 27924 14297 27939
rect 14331 27924 14361 27958
rect 13968 27901 14361 27924
rect 13968 27867 14122 27901
rect 14156 27890 14361 27901
rect 14156 27867 14297 27890
rect 13968 27856 14297 27867
rect 14331 27856 14361 27890
rect 13968 27829 14361 27856
rect 13968 27795 14122 27829
rect 14156 27822 14361 27829
rect 14156 27795 14297 27822
rect 13968 27788 14297 27795
rect 14331 27788 14361 27822
rect 13968 27757 14361 27788
rect 13968 27723 14122 27757
rect 14156 27754 14361 27757
rect 14156 27723 14297 27754
rect 13968 27720 14297 27723
rect 14331 27720 14361 27754
rect 13968 27686 14361 27720
rect 13968 27685 14297 27686
rect 13968 27651 14122 27685
rect 14156 27652 14297 27685
rect 14331 27652 14361 27686
rect 14156 27651 14361 27652
rect 13968 27618 14361 27651
rect 13968 27613 14297 27618
rect 13968 27579 14122 27613
rect 14156 27584 14297 27613
rect 14331 27584 14361 27618
rect 14156 27579 14361 27584
rect 13968 27550 14361 27579
rect 13968 27541 14297 27550
rect 13968 27507 14122 27541
rect 14156 27516 14297 27541
rect 14331 27516 14361 27550
rect 14156 27507 14361 27516
rect 13968 27482 14361 27507
rect 13968 27469 14297 27482
rect 13968 27435 14122 27469
rect 14156 27448 14297 27469
rect 14331 27448 14361 27482
rect 14156 27435 14361 27448
rect 13968 27414 14361 27435
rect 13968 27397 14297 27414
rect 13968 27363 14122 27397
rect 14156 27380 14297 27397
rect 14331 27380 14361 27414
rect 14156 27363 14361 27380
rect 13968 27346 14361 27363
rect 13968 27325 14297 27346
rect 13968 27291 14122 27325
rect 14156 27312 14297 27325
rect 14331 27312 14361 27346
rect 14156 27291 14361 27312
rect 13968 27278 14361 27291
rect 13968 27253 14297 27278
rect 13968 27219 14122 27253
rect 14156 27244 14297 27253
rect 14331 27244 14361 27278
rect 14156 27219 14361 27244
rect 13968 27210 14361 27219
rect 13968 27181 14297 27210
rect 13968 27147 14122 27181
rect 14156 27176 14297 27181
rect 14331 27176 14361 27210
rect 14156 27147 14361 27176
rect 13968 27142 14361 27147
rect 13968 27109 14297 27142
rect 13968 27075 14122 27109
rect 14156 27108 14297 27109
rect 14331 27108 14361 27142
rect 14156 27075 14361 27108
rect 13968 27074 14361 27075
rect 13968 27040 14297 27074
rect 14331 27040 14361 27074
rect 13968 27037 14361 27040
rect 13968 27003 14122 27037
rect 14156 27006 14361 27037
rect 14156 27003 14297 27006
rect 13968 26972 14297 27003
rect 14331 26972 14361 27006
rect 13968 26965 14361 26972
rect 13968 26931 14122 26965
rect 14156 26938 14361 26965
rect 14156 26931 14297 26938
rect 13968 26904 14297 26931
rect 14331 26904 14361 26938
rect 13968 26893 14361 26904
rect 13968 26859 14122 26893
rect 14156 26870 14361 26893
rect 14156 26859 14297 26870
rect 13968 26836 14297 26859
rect 14331 26836 14361 26870
rect 13968 26821 14361 26836
rect 13968 26787 14122 26821
rect 14156 26802 14361 26821
rect 14156 26787 14297 26802
rect 13968 26768 14297 26787
rect 14331 26768 14361 26802
rect 13968 26749 14361 26768
rect 13968 26715 14122 26749
rect 14156 26734 14361 26749
rect 14156 26715 14297 26734
rect 13968 26700 14297 26715
rect 14331 26700 14361 26734
rect 13968 26677 14361 26700
rect 13968 26643 14122 26677
rect 14156 26666 14361 26677
rect 14156 26643 14297 26666
rect 13968 26632 14297 26643
rect 14331 26632 14361 26666
rect 13968 26605 14361 26632
rect 13968 26571 14122 26605
rect 14156 26598 14361 26605
rect 14156 26571 14297 26598
rect 13968 26564 14297 26571
rect 14331 26564 14361 26598
rect 13968 26533 14361 26564
rect 13968 26499 14122 26533
rect 14156 26530 14361 26533
rect 14156 26499 14297 26530
rect 13968 26496 14297 26499
rect 14331 26496 14361 26530
rect 13968 26462 14361 26496
rect 13968 26461 14297 26462
rect 13968 26427 14122 26461
rect 14156 26428 14297 26461
rect 14331 26428 14361 26462
rect 14156 26427 14361 26428
rect 13968 26394 14361 26427
rect 13968 26389 14297 26394
rect 13968 26355 14122 26389
rect 14156 26360 14297 26389
rect 14331 26360 14361 26394
rect 14156 26355 14361 26360
rect 13968 26326 14361 26355
rect 13968 26317 14297 26326
rect 13968 26283 14122 26317
rect 14156 26292 14297 26317
rect 14331 26292 14361 26326
rect 14156 26283 14361 26292
rect 13968 26258 14361 26283
rect 13968 26245 14297 26258
rect 13968 26211 14122 26245
rect 14156 26224 14297 26245
rect 14331 26224 14361 26258
rect 14156 26211 14361 26224
rect 13968 26190 14361 26211
rect 13968 26173 14297 26190
rect 13968 26139 14122 26173
rect 14156 26156 14297 26173
rect 14331 26156 14361 26190
rect 14156 26139 14361 26156
rect 13968 26122 14361 26139
rect 13968 26101 14297 26122
rect 13968 26067 14122 26101
rect 14156 26088 14297 26101
rect 14331 26088 14361 26122
rect 14156 26067 14361 26088
rect 13968 26054 14361 26067
rect 13968 26029 14297 26054
rect 13968 25995 14122 26029
rect 14156 26020 14297 26029
rect 14331 26020 14361 26054
rect 14156 25995 14361 26020
rect 13968 25986 14361 25995
rect 13968 25957 14297 25986
rect 13968 25923 14122 25957
rect 14156 25952 14297 25957
rect 14331 25952 14361 25986
rect 14156 25923 14361 25952
rect 13968 25918 14361 25923
rect 13968 25885 14297 25918
rect 13968 25851 14122 25885
rect 14156 25884 14297 25885
rect 14331 25884 14361 25918
rect 14156 25851 14361 25884
rect 13968 25850 14361 25851
rect 13968 25816 14297 25850
rect 14331 25816 14361 25850
rect 13968 25813 14361 25816
rect 13968 25779 14122 25813
rect 14156 25782 14361 25813
rect 14156 25779 14297 25782
rect 13968 25748 14297 25779
rect 14331 25748 14361 25782
rect 13968 25741 14361 25748
rect 13968 25707 14122 25741
rect 14156 25714 14361 25741
rect 14156 25707 14297 25714
rect 13968 25680 14297 25707
rect 14331 25680 14361 25714
rect 13968 25669 14361 25680
rect 13968 25635 14122 25669
rect 14156 25646 14361 25669
rect 14156 25635 14297 25646
rect 13968 25612 14297 25635
rect 14331 25612 14361 25646
rect 13968 25597 14361 25612
rect 13968 25563 14122 25597
rect 14156 25578 14361 25597
rect 14156 25563 14297 25578
rect 13968 25544 14297 25563
rect 14331 25544 14361 25578
rect 13968 25525 14361 25544
rect 13968 25491 14122 25525
rect 14156 25510 14361 25525
rect 14156 25491 14297 25510
rect 13968 25476 14297 25491
rect 14331 25476 14361 25510
rect 13968 25453 14361 25476
rect 13968 25419 14122 25453
rect 14156 25442 14361 25453
rect 14156 25419 14297 25442
rect 13968 25408 14297 25419
rect 14331 25408 14361 25442
rect 13968 25381 14361 25408
rect 13968 25347 14122 25381
rect 14156 25374 14361 25381
rect 14156 25347 14297 25374
rect 13968 25340 14297 25347
rect 14331 25340 14361 25374
rect 13968 25309 14361 25340
rect 13968 25275 14122 25309
rect 14156 25306 14361 25309
rect 14156 25275 14297 25306
rect 13968 25272 14297 25275
rect 14331 25272 14361 25306
rect 13968 25238 14361 25272
rect 13968 25237 14297 25238
rect 13968 25203 14122 25237
rect 14156 25204 14297 25237
rect 14331 25204 14361 25238
rect 14156 25203 14361 25204
rect 13968 25170 14361 25203
rect 13968 25165 14297 25170
rect 13968 25131 14122 25165
rect 14156 25136 14297 25165
rect 14331 25136 14361 25170
rect 14156 25131 14361 25136
rect 13968 25102 14361 25131
rect 13968 25093 14297 25102
rect 13968 25059 14122 25093
rect 14156 25068 14297 25093
rect 14331 25068 14361 25102
rect 14156 25059 14361 25068
rect 13968 25034 14361 25059
rect 13968 25021 14297 25034
rect 13968 24987 14122 25021
rect 14156 25000 14297 25021
rect 14331 25000 14361 25034
rect 14156 24987 14361 25000
rect 13968 24966 14361 24987
rect 13968 24949 14297 24966
rect 13968 24915 14122 24949
rect 14156 24932 14297 24949
rect 14331 24932 14361 24966
rect 14156 24915 14361 24932
rect 13968 24898 14361 24915
rect 13968 24877 14297 24898
rect 13968 24843 14122 24877
rect 14156 24864 14297 24877
rect 14331 24864 14361 24898
rect 14156 24843 14361 24864
rect 13968 24830 14361 24843
rect 13968 24805 14297 24830
rect 13968 24771 14122 24805
rect 14156 24796 14297 24805
rect 14331 24796 14361 24830
rect 14156 24771 14361 24796
rect 13968 24762 14361 24771
rect 13968 24733 14297 24762
rect 13968 24699 14122 24733
rect 14156 24728 14297 24733
rect 14331 24728 14361 24762
rect 14156 24699 14361 24728
rect 13968 24694 14361 24699
rect 13968 24661 14297 24694
rect 13968 24627 14122 24661
rect 14156 24660 14297 24661
rect 14331 24660 14361 24694
rect 14156 24627 14361 24660
rect 13968 24626 14361 24627
rect 13968 24592 14297 24626
rect 14331 24592 14361 24626
rect 13968 24589 14361 24592
rect 13968 24555 14122 24589
rect 14156 24558 14361 24589
rect 14156 24555 14297 24558
rect 13968 24524 14297 24555
rect 14331 24524 14361 24558
rect 13968 24517 14361 24524
rect 13968 24483 14122 24517
rect 14156 24490 14361 24517
rect 14156 24483 14297 24490
rect 13968 24456 14297 24483
rect 14331 24456 14361 24490
rect 13968 24445 14361 24456
rect 13968 24411 14122 24445
rect 14156 24422 14361 24445
rect 14156 24411 14297 24422
rect 13968 24388 14297 24411
rect 14331 24388 14361 24422
rect 13968 24373 14361 24388
rect 13968 24339 14122 24373
rect 14156 24354 14361 24373
rect 14156 24339 14297 24354
rect 13968 24320 14297 24339
rect 14331 24320 14361 24354
rect 13968 24301 14361 24320
rect 13968 24267 14122 24301
rect 14156 24286 14361 24301
rect 14156 24267 14297 24286
rect 13968 24252 14297 24267
rect 14331 24252 14361 24286
rect 13968 24229 14361 24252
rect 13968 24195 14122 24229
rect 14156 24218 14361 24229
rect 14156 24195 14297 24218
rect 13968 24184 14297 24195
rect 14331 24184 14361 24218
rect 13968 24157 14361 24184
rect 13968 24123 14122 24157
rect 14156 24150 14361 24157
rect 14156 24123 14297 24150
rect 13968 24116 14297 24123
rect 14331 24116 14361 24150
rect 13968 24085 14361 24116
rect 13968 24051 14122 24085
rect 14156 24082 14361 24085
rect 14156 24051 14297 24082
rect 13968 24048 14297 24051
rect 14331 24048 14361 24082
rect 13968 24014 14361 24048
rect 13968 24013 14297 24014
rect 13968 23979 14122 24013
rect 14156 23980 14297 24013
rect 14331 23980 14361 24014
rect 14156 23979 14361 23980
rect 13968 23946 14361 23979
rect 13968 23941 14297 23946
rect 13968 23907 14122 23941
rect 14156 23912 14297 23941
rect 14331 23912 14361 23946
rect 14156 23907 14361 23912
rect 13968 23878 14361 23907
rect 13968 23869 14297 23878
rect 13968 23835 14122 23869
rect 14156 23844 14297 23869
rect 14331 23844 14361 23878
rect 14156 23835 14361 23844
rect 13968 23810 14361 23835
rect 13968 23797 14297 23810
rect 13968 23763 14122 23797
rect 14156 23776 14297 23797
rect 14331 23776 14361 23810
rect 14156 23763 14361 23776
rect 13968 23742 14361 23763
rect 13968 23725 14297 23742
rect 13968 23691 14122 23725
rect 14156 23708 14297 23725
rect 14331 23708 14361 23742
rect 14156 23691 14361 23708
rect 13968 23674 14361 23691
rect 13968 23653 14297 23674
rect 13968 23619 14122 23653
rect 14156 23640 14297 23653
rect 14331 23640 14361 23674
rect 14156 23619 14361 23640
rect 13968 23606 14361 23619
rect 13968 23581 14297 23606
rect 13968 23547 14122 23581
rect 14156 23572 14297 23581
rect 14331 23572 14361 23606
rect 14156 23547 14361 23572
rect 13968 23538 14361 23547
rect 13968 23509 14297 23538
rect 13968 23475 14122 23509
rect 14156 23504 14297 23509
rect 14331 23504 14361 23538
rect 14156 23475 14361 23504
rect 13968 23470 14361 23475
rect 13968 23437 14297 23470
rect 13968 23403 14122 23437
rect 14156 23436 14297 23437
rect 14331 23436 14361 23470
rect 14156 23403 14361 23436
rect 13968 23402 14361 23403
rect 13968 23368 14297 23402
rect 14331 23368 14361 23402
rect 13968 23365 14361 23368
rect 13968 23331 14122 23365
rect 14156 23334 14361 23365
rect 14156 23331 14297 23334
rect 13968 23300 14297 23331
rect 14331 23300 14361 23334
rect 13968 23293 14361 23300
rect 13968 23259 14122 23293
rect 14156 23266 14361 23293
rect 14156 23259 14297 23266
rect 13968 23232 14297 23259
rect 14331 23232 14361 23266
rect 13968 23221 14361 23232
rect 13968 23187 14122 23221
rect 14156 23198 14361 23221
rect 14156 23187 14297 23198
rect 13968 23164 14297 23187
rect 14331 23164 14361 23198
rect 13968 23149 14361 23164
rect 13968 23115 14122 23149
rect 14156 23130 14361 23149
rect 14156 23115 14297 23130
rect 13968 23096 14297 23115
rect 14331 23096 14361 23130
rect 13968 23077 14361 23096
rect 13968 23043 14122 23077
rect 14156 23062 14361 23077
rect 14156 23043 14297 23062
rect 13968 23028 14297 23043
rect 14331 23028 14361 23062
rect 13968 23005 14361 23028
rect 13968 22971 14122 23005
rect 14156 22994 14361 23005
rect 14156 22971 14297 22994
rect 13968 22960 14297 22971
rect 14331 22960 14361 22994
rect 13968 22933 14361 22960
rect 13968 22899 14122 22933
rect 14156 22926 14361 22933
rect 14156 22899 14297 22926
rect 13968 22892 14297 22899
rect 14331 22892 14361 22926
rect 13968 22861 14361 22892
rect 13968 22827 14122 22861
rect 14156 22858 14361 22861
rect 14156 22827 14297 22858
rect 13968 22824 14297 22827
rect 14331 22824 14361 22858
rect 13968 22790 14361 22824
rect 13968 22789 14297 22790
rect 13968 22755 14122 22789
rect 14156 22756 14297 22789
rect 14331 22756 14361 22790
rect 14156 22755 14361 22756
rect 13968 22722 14361 22755
rect 13968 22717 14297 22722
rect 13968 22683 14122 22717
rect 14156 22688 14297 22717
rect 14331 22688 14361 22722
rect 14156 22683 14361 22688
rect 13968 22654 14361 22683
rect 13968 22645 14297 22654
rect 13968 22611 14122 22645
rect 14156 22620 14297 22645
rect 14331 22620 14361 22654
rect 14156 22611 14361 22620
rect 13968 22586 14361 22611
rect 13968 22573 14297 22586
rect 13968 22539 14122 22573
rect 14156 22552 14297 22573
rect 14331 22552 14361 22586
rect 14156 22539 14361 22552
rect 13968 22518 14361 22539
rect 13968 22501 14297 22518
rect 13968 22467 14122 22501
rect 14156 22484 14297 22501
rect 14331 22484 14361 22518
rect 14156 22467 14361 22484
rect 13968 22450 14361 22467
rect 13968 22429 14297 22450
rect 13968 22395 14122 22429
rect 14156 22416 14297 22429
rect 14331 22416 14361 22450
rect 14156 22395 14361 22416
rect 13968 22382 14361 22395
rect 13968 22357 14297 22382
rect 13968 22323 14122 22357
rect 14156 22348 14297 22357
rect 14331 22348 14361 22382
rect 14156 22323 14361 22348
rect 13968 22314 14361 22323
rect 13968 22285 14297 22314
rect 13968 22251 14122 22285
rect 14156 22280 14297 22285
rect 14331 22280 14361 22314
rect 14156 22251 14361 22280
rect 13968 22246 14361 22251
rect 13968 22213 14297 22246
rect 13968 22179 14122 22213
rect 14156 22212 14297 22213
rect 14331 22212 14361 22246
rect 14156 22179 14361 22212
rect 13968 22178 14361 22179
rect 13968 22144 14297 22178
rect 14331 22144 14361 22178
rect 13968 22141 14361 22144
rect 13968 22107 14122 22141
rect 14156 22110 14361 22141
rect 14156 22107 14297 22110
rect 13968 22076 14297 22107
rect 14331 22076 14361 22110
rect 13968 22069 14361 22076
rect 13968 22035 14122 22069
rect 14156 22042 14361 22069
rect 14156 22035 14297 22042
rect 13968 22008 14297 22035
rect 14331 22008 14361 22042
rect 13968 21997 14361 22008
rect 13968 21963 14122 21997
rect 14156 21974 14361 21997
rect 14156 21963 14297 21974
rect 13968 21940 14297 21963
rect 14331 21940 14361 21974
rect 13968 21925 14361 21940
rect 13968 21891 14122 21925
rect 14156 21906 14361 21925
rect 14156 21891 14297 21906
rect 13968 21872 14297 21891
rect 14331 21872 14361 21906
rect 13968 21853 14361 21872
rect 13968 21819 14122 21853
rect 14156 21838 14361 21853
rect 14156 21819 14297 21838
rect 13968 21804 14297 21819
rect 14331 21804 14361 21838
rect 13968 21781 14361 21804
rect 13968 21747 14122 21781
rect 14156 21770 14361 21781
rect 14156 21747 14297 21770
rect 13968 21736 14297 21747
rect 14331 21736 14361 21770
rect 13968 21709 14361 21736
rect 13968 21675 14122 21709
rect 14156 21702 14361 21709
rect 14156 21675 14297 21702
rect 13968 21668 14297 21675
rect 14331 21668 14361 21702
rect 13968 21637 14361 21668
rect 13968 21603 14122 21637
rect 14156 21634 14361 21637
rect 14156 21603 14297 21634
rect 13968 21600 14297 21603
rect 14331 21600 14361 21634
rect 13968 21566 14361 21600
rect 13968 21565 14297 21566
rect 13968 21531 14122 21565
rect 14156 21532 14297 21565
rect 14331 21532 14361 21566
rect 14156 21531 14361 21532
rect 13968 21498 14361 21531
rect 13968 21493 14297 21498
rect 13968 21459 14122 21493
rect 14156 21464 14297 21493
rect 14331 21464 14361 21498
rect 14156 21459 14361 21464
rect 13968 21430 14361 21459
rect 13968 21421 14297 21430
rect 13968 21387 14122 21421
rect 14156 21396 14297 21421
rect 14331 21396 14361 21430
rect 14156 21387 14361 21396
rect 13968 21362 14361 21387
rect 13968 21349 14297 21362
rect 13968 21315 14122 21349
rect 14156 21328 14297 21349
rect 14331 21328 14361 21362
rect 14156 21315 14361 21328
rect 13968 21294 14361 21315
rect 13968 21277 14297 21294
rect 13968 21243 14122 21277
rect 14156 21260 14297 21277
rect 14331 21260 14361 21294
rect 14156 21243 14361 21260
rect 13968 21226 14361 21243
rect 13968 21205 14297 21226
rect 13968 21171 14122 21205
rect 14156 21192 14297 21205
rect 14331 21192 14361 21226
rect 14156 21171 14361 21192
rect 13968 21158 14361 21171
rect 13968 21133 14297 21158
rect 13968 21099 14122 21133
rect 14156 21124 14297 21133
rect 14331 21124 14361 21158
rect 14156 21099 14361 21124
rect 13968 21090 14361 21099
rect 13968 21061 14297 21090
rect 13968 21027 14122 21061
rect 14156 21056 14297 21061
rect 14331 21056 14361 21090
rect 14156 21027 14361 21056
rect 13968 21022 14361 21027
rect 13968 20989 14297 21022
rect 13968 20955 14122 20989
rect 14156 20988 14297 20989
rect 14331 20988 14361 21022
rect 14156 20955 14361 20988
rect 13968 20954 14361 20955
rect 13968 20920 14297 20954
rect 14331 20920 14361 20954
rect 13968 20917 14361 20920
rect 13968 20883 14122 20917
rect 14156 20886 14361 20917
rect 14156 20883 14297 20886
rect 13968 20852 14297 20883
rect 14331 20852 14361 20886
rect 13968 20845 14361 20852
rect 13968 20811 14122 20845
rect 14156 20818 14361 20845
rect 14156 20811 14297 20818
rect 13968 20784 14297 20811
rect 14331 20784 14361 20818
rect 13968 20773 14361 20784
rect 13968 20739 14122 20773
rect 14156 20750 14361 20773
rect 14156 20739 14297 20750
rect 13968 20716 14297 20739
rect 14331 20716 14361 20750
rect 13968 20701 14361 20716
rect 13968 20667 14122 20701
rect 14156 20682 14361 20701
rect 14156 20667 14297 20682
rect 13968 20648 14297 20667
rect 14331 20648 14361 20682
rect 13968 20629 14361 20648
rect 13968 20595 14122 20629
rect 14156 20614 14361 20629
rect 14156 20595 14297 20614
rect 13968 20580 14297 20595
rect 14331 20580 14361 20614
rect 13968 20557 14361 20580
rect 13968 20523 14122 20557
rect 14156 20546 14361 20557
rect 14156 20523 14297 20546
rect 13968 20512 14297 20523
rect 14331 20512 14361 20546
rect 13968 20485 14361 20512
rect 13968 20451 14122 20485
rect 14156 20478 14361 20485
rect 14156 20451 14297 20478
rect 13968 20444 14297 20451
rect 14331 20444 14361 20478
rect 13968 20413 14361 20444
rect 13968 20379 14122 20413
rect 14156 20410 14361 20413
rect 14156 20379 14297 20410
rect 13968 20376 14297 20379
rect 14331 20376 14361 20410
rect 13968 20342 14361 20376
rect 13968 20341 14297 20342
rect 13968 20307 14122 20341
rect 14156 20308 14297 20341
rect 14331 20308 14361 20342
rect 14156 20307 14361 20308
rect 13968 20274 14361 20307
rect 13968 20269 14297 20274
rect 13968 20235 14122 20269
rect 14156 20240 14297 20269
rect 14331 20240 14361 20274
rect 14156 20235 14361 20240
rect 13968 20206 14361 20235
rect 13968 20197 14297 20206
rect 13968 20163 14122 20197
rect 14156 20172 14297 20197
rect 14331 20172 14361 20206
rect 14156 20163 14361 20172
rect 13968 20138 14361 20163
rect 13968 20125 14297 20138
rect 13968 20091 14122 20125
rect 14156 20104 14297 20125
rect 14331 20104 14361 20138
rect 14156 20091 14361 20104
rect 13968 20070 14361 20091
rect 13968 20053 14297 20070
rect 13968 20019 14122 20053
rect 14156 20036 14297 20053
rect 14331 20036 14361 20070
rect 14156 20019 14361 20036
rect 13968 20002 14361 20019
rect 13968 19981 14297 20002
rect 13968 19947 14122 19981
rect 14156 19968 14297 19981
rect 14331 19968 14361 20002
rect 14156 19947 14361 19968
rect 13968 19934 14361 19947
rect 13968 19909 14297 19934
rect 13968 19875 14122 19909
rect 14156 19900 14297 19909
rect 14331 19900 14361 19934
rect 14156 19875 14361 19900
rect 13968 19866 14361 19875
rect 13968 19837 14297 19866
rect 13968 19803 14122 19837
rect 14156 19832 14297 19837
rect 14331 19832 14361 19866
rect 14156 19803 14361 19832
rect 13968 19798 14361 19803
rect 13968 19765 14297 19798
rect 13968 19731 14122 19765
rect 14156 19764 14297 19765
rect 14331 19764 14361 19798
rect 14156 19731 14361 19764
rect 13968 19730 14361 19731
rect 13968 19696 14297 19730
rect 14331 19696 14361 19730
rect 13968 19693 14361 19696
rect 13968 19659 14122 19693
rect 14156 19662 14361 19693
rect 14156 19659 14297 19662
rect 13968 19628 14297 19659
rect 14331 19628 14361 19662
rect 13968 19621 14361 19628
rect 13968 19587 14122 19621
rect 14156 19594 14361 19621
rect 14156 19587 14297 19594
rect 13968 19560 14297 19587
rect 14331 19560 14361 19594
rect 13968 19549 14361 19560
rect 13968 19515 14122 19549
rect 14156 19526 14361 19549
rect 14156 19515 14297 19526
rect 13968 19492 14297 19515
rect 14331 19492 14361 19526
rect 13968 19477 14361 19492
rect 13968 19443 14122 19477
rect 14156 19458 14361 19477
rect 14156 19443 14297 19458
rect 13968 19424 14297 19443
rect 14331 19424 14361 19458
rect 13968 19405 14361 19424
rect 13968 19371 14122 19405
rect 14156 19390 14361 19405
rect 14156 19371 14297 19390
rect 13968 19356 14297 19371
rect 14331 19356 14361 19390
rect 13968 19333 14361 19356
rect 13968 19299 14122 19333
rect 14156 19322 14361 19333
rect 14156 19299 14297 19322
rect 13968 19288 14297 19299
rect 14331 19288 14361 19322
rect 13968 19261 14361 19288
rect 13968 19227 14122 19261
rect 14156 19254 14361 19261
rect 14156 19227 14297 19254
rect 13968 19220 14297 19227
rect 14331 19220 14361 19254
rect 13968 19189 14361 19220
rect 13968 19155 14122 19189
rect 14156 19186 14361 19189
rect 14156 19155 14297 19186
rect 13968 19152 14297 19155
rect 14331 19152 14361 19186
rect 13968 19118 14361 19152
rect 13968 19117 14297 19118
rect 13968 19083 14122 19117
rect 14156 19084 14297 19117
rect 14331 19084 14361 19118
rect 14156 19083 14361 19084
rect 13968 19050 14361 19083
rect 13968 19045 14297 19050
rect 13968 19011 14122 19045
rect 14156 19016 14297 19045
rect 14331 19016 14361 19050
rect 14156 19011 14361 19016
rect 13968 18982 14361 19011
rect 13968 18973 14297 18982
rect 13968 18939 14122 18973
rect 14156 18948 14297 18973
rect 14331 18948 14361 18982
rect 14156 18939 14361 18948
rect 13968 18914 14361 18939
rect 13968 18901 14297 18914
rect 13968 18867 14122 18901
rect 14156 18880 14297 18901
rect 14331 18880 14361 18914
rect 14156 18867 14361 18880
rect 13968 18846 14361 18867
rect 13968 18829 14297 18846
rect 13968 18795 14122 18829
rect 14156 18812 14297 18829
rect 14331 18812 14361 18846
rect 14156 18795 14361 18812
rect 13968 18778 14361 18795
rect 13968 18757 14297 18778
rect 13968 18723 14122 18757
rect 14156 18744 14297 18757
rect 14331 18744 14361 18778
rect 14156 18723 14361 18744
rect 13968 18710 14361 18723
rect 13968 18685 14297 18710
rect 13968 18651 14122 18685
rect 14156 18676 14297 18685
rect 14331 18676 14361 18710
rect 14156 18651 14361 18676
rect 13968 18642 14361 18651
rect 13968 18613 14297 18642
rect 13968 18579 14122 18613
rect 14156 18608 14297 18613
rect 14331 18608 14361 18642
rect 14156 18579 14361 18608
rect 13968 18574 14361 18579
rect 13968 18541 14297 18574
rect 13968 18507 14122 18541
rect 14156 18540 14297 18541
rect 14331 18540 14361 18574
rect 14156 18507 14361 18540
rect 13968 18506 14361 18507
rect 13968 18472 14297 18506
rect 14331 18472 14361 18506
rect 13968 18469 14361 18472
rect 13968 18435 14122 18469
rect 14156 18438 14361 18469
rect 14156 18435 14297 18438
rect 13968 18404 14297 18435
rect 14331 18404 14361 18438
rect 13968 18397 14361 18404
rect 13968 18363 14122 18397
rect 14156 18370 14361 18397
rect 14156 18363 14297 18370
rect 13968 18336 14297 18363
rect 14331 18336 14361 18370
rect 13968 18325 14361 18336
rect 13968 18291 14122 18325
rect 14156 18302 14361 18325
rect 14156 18291 14297 18302
rect 13968 18268 14297 18291
rect 14331 18268 14361 18302
rect 13968 18253 14361 18268
rect 13968 18219 14122 18253
rect 14156 18234 14361 18253
rect 14156 18219 14297 18234
rect 13968 18200 14297 18219
rect 14331 18200 14361 18234
rect 13968 18181 14361 18200
rect 13968 18147 14122 18181
rect 14156 18166 14361 18181
rect 14156 18147 14297 18166
rect 13968 18132 14297 18147
rect 14331 18132 14361 18166
rect 13968 18109 14361 18132
rect 13968 18075 14122 18109
rect 14156 18098 14361 18109
rect 14156 18075 14297 18098
rect 13968 18064 14297 18075
rect 14331 18064 14361 18098
rect 13968 18037 14361 18064
rect 13968 18003 14122 18037
rect 14156 18030 14361 18037
rect 14156 18003 14297 18030
rect 13968 17996 14297 18003
rect 14331 17996 14361 18030
rect 13968 17965 14361 17996
rect 13968 17931 14122 17965
rect 14156 17962 14361 17965
rect 14156 17931 14297 17962
rect 13968 17928 14297 17931
rect 14331 17928 14361 17962
rect 13968 17894 14361 17928
rect 13968 17893 14297 17894
rect 13968 17859 14122 17893
rect 14156 17860 14297 17893
rect 14331 17860 14361 17894
rect 14156 17859 14361 17860
rect 13968 17826 14361 17859
rect 13968 17821 14297 17826
rect 13968 17787 14122 17821
rect 14156 17792 14297 17821
rect 14331 17792 14361 17826
rect 14156 17787 14361 17792
rect 13968 17758 14361 17787
rect 13968 17749 14297 17758
rect 13968 17715 14122 17749
rect 14156 17724 14297 17749
rect 14331 17724 14361 17758
rect 14156 17715 14361 17724
rect 13968 17690 14361 17715
rect 13968 17677 14297 17690
rect 13968 17643 14122 17677
rect 14156 17656 14297 17677
rect 14331 17656 14361 17690
rect 14156 17643 14361 17656
rect 13968 17622 14361 17643
rect 13968 17605 14297 17622
rect 13968 17571 14122 17605
rect 14156 17588 14297 17605
rect 14331 17588 14361 17622
rect 14156 17571 14361 17588
rect 13968 17554 14361 17571
rect 13968 17533 14297 17554
rect 13968 17499 14122 17533
rect 14156 17520 14297 17533
rect 14331 17520 14361 17554
rect 14156 17499 14361 17520
rect 13968 17486 14361 17499
rect 13968 17461 14297 17486
rect 13968 17427 14122 17461
rect 14156 17452 14297 17461
rect 14331 17452 14361 17486
rect 14156 17427 14361 17452
rect 13968 17418 14361 17427
rect 13968 17389 14297 17418
rect 13968 17355 14122 17389
rect 14156 17384 14297 17389
rect 14331 17384 14361 17418
rect 14156 17355 14361 17384
rect 13968 17350 14361 17355
rect 13968 17317 14297 17350
rect 13968 17283 14122 17317
rect 14156 17316 14297 17317
rect 14331 17316 14361 17350
rect 14156 17283 14361 17316
rect 13968 17282 14361 17283
rect 13968 17248 14297 17282
rect 14331 17248 14361 17282
rect 13968 17245 14361 17248
rect 13968 17211 14122 17245
rect 14156 17214 14361 17245
rect 14156 17211 14297 17214
rect 13968 17180 14297 17211
rect 14331 17180 14361 17214
rect 13968 17173 14361 17180
rect 13968 17139 14122 17173
rect 14156 17146 14361 17173
rect 14156 17139 14297 17146
rect 13968 17112 14297 17139
rect 14331 17112 14361 17146
rect 13968 17101 14361 17112
rect 13968 17067 14122 17101
rect 14156 17078 14361 17101
rect 14156 17067 14297 17078
rect 13968 17044 14297 17067
rect 14331 17044 14361 17078
rect 13968 17029 14361 17044
rect 13968 16995 14122 17029
rect 14156 17010 14361 17029
rect 14156 16995 14297 17010
rect 13968 16976 14297 16995
rect 14331 16976 14361 17010
rect 13968 16957 14361 16976
rect 13968 16923 14122 16957
rect 14156 16942 14361 16957
rect 14156 16923 14297 16942
rect 13968 16908 14297 16923
rect 14331 16908 14361 16942
rect 13968 16885 14361 16908
rect 13968 16851 14122 16885
rect 14156 16874 14361 16885
rect 14156 16851 14297 16874
rect 13968 16840 14297 16851
rect 14331 16840 14361 16874
rect 13968 16813 14361 16840
rect 13968 16779 14122 16813
rect 14156 16806 14361 16813
rect 14156 16779 14297 16806
rect 13968 16772 14297 16779
rect 14331 16772 14361 16806
rect 13968 16741 14361 16772
rect 13968 16707 14122 16741
rect 14156 16738 14361 16741
rect 14156 16707 14297 16738
rect 13968 16704 14297 16707
rect 14331 16704 14361 16738
rect 13968 16670 14361 16704
rect 13968 16669 14297 16670
rect 13968 16635 14122 16669
rect 14156 16636 14297 16669
rect 14331 16636 14361 16670
rect 14156 16635 14361 16636
rect 13968 16602 14361 16635
rect 13968 16597 14297 16602
rect 13968 16563 14122 16597
rect 14156 16568 14297 16597
rect 14331 16568 14361 16602
rect 14156 16563 14361 16568
rect 13968 16534 14361 16563
rect 13968 16525 14297 16534
rect 13968 16491 14122 16525
rect 14156 16500 14297 16525
rect 14331 16500 14361 16534
rect 14156 16491 14361 16500
rect 13968 16466 14361 16491
rect 13968 16453 14297 16466
rect 13968 16419 14122 16453
rect 14156 16432 14297 16453
rect 14331 16432 14361 16466
rect 14156 16419 14361 16432
rect 13968 16398 14361 16419
rect 13968 16381 14297 16398
rect 13968 16347 14122 16381
rect 14156 16364 14297 16381
rect 14331 16364 14361 16398
rect 14156 16347 14361 16364
rect 13968 16330 14361 16347
rect 13968 16309 14297 16330
rect 13968 16275 14122 16309
rect 14156 16296 14297 16309
rect 14331 16296 14361 16330
rect 14156 16275 14361 16296
rect 13968 16262 14361 16275
rect 13968 16237 14297 16262
rect 13968 16203 14122 16237
rect 14156 16228 14297 16237
rect 14331 16228 14361 16262
rect 14156 16203 14361 16228
rect 13968 16194 14361 16203
rect 13968 16165 14297 16194
rect 13968 16131 14122 16165
rect 14156 16160 14297 16165
rect 14331 16160 14361 16194
rect 14156 16131 14361 16160
rect 13968 16126 14361 16131
rect 13968 16093 14297 16126
rect 13968 16059 14122 16093
rect 14156 16092 14297 16093
rect 14331 16092 14361 16126
rect 14156 16059 14361 16092
rect 13968 16058 14361 16059
rect 13968 16024 14297 16058
rect 14331 16024 14361 16058
rect 13968 16021 14361 16024
rect 13968 15987 14122 16021
rect 14156 15990 14361 16021
rect 14156 15987 14297 15990
rect 13968 15956 14297 15987
rect 14331 15956 14361 15990
rect 13968 15949 14361 15956
rect 13968 15915 14122 15949
rect 14156 15922 14361 15949
rect 14156 15915 14297 15922
rect 13968 15888 14297 15915
rect 14331 15888 14361 15922
rect 13968 15877 14361 15888
rect 13968 15843 14122 15877
rect 14156 15854 14361 15877
rect 14156 15843 14297 15854
rect 13968 15820 14297 15843
rect 14331 15820 14361 15854
rect 13968 15805 14361 15820
rect 13968 15771 14122 15805
rect 14156 15786 14361 15805
rect 14156 15771 14297 15786
rect 13968 15752 14297 15771
rect 14331 15752 14361 15786
rect 13968 15733 14361 15752
rect 13968 15699 14122 15733
rect 14156 15718 14361 15733
rect 14156 15699 14297 15718
rect 13968 15684 14297 15699
rect 14331 15684 14361 15718
rect 13968 15661 14361 15684
rect 13968 15627 14122 15661
rect 14156 15650 14361 15661
rect 14156 15627 14297 15650
rect 13968 15616 14297 15627
rect 14331 15616 14361 15650
rect 13968 15589 14361 15616
rect 13968 15555 14122 15589
rect 14156 15582 14361 15589
rect 14156 15555 14297 15582
rect 13968 15548 14297 15555
rect 14331 15548 14361 15582
rect 13968 15517 14361 15548
rect 13968 15483 14122 15517
rect 14156 15514 14361 15517
rect 14156 15483 14297 15514
rect 13968 15480 14297 15483
rect 14331 15480 14361 15514
rect 13968 15446 14361 15480
rect 13968 15445 14297 15446
rect 13968 15411 14122 15445
rect 14156 15412 14297 15445
rect 14331 15412 14361 15446
rect 14156 15411 14361 15412
rect 13968 15378 14361 15411
rect 13968 15373 14297 15378
rect 13968 15339 14122 15373
rect 14156 15344 14297 15373
rect 14331 15344 14361 15378
rect 14156 15339 14361 15344
rect 13968 15310 14361 15339
rect 13968 15301 14297 15310
rect 13968 15267 14122 15301
rect 14156 15276 14297 15301
rect 14331 15276 14361 15310
rect 14156 15267 14361 15276
rect 13968 15242 14361 15267
rect 13968 15229 14297 15242
rect 603 15140 632 15174
rect 666 15164 1026 15174
rect 666 15140 807 15164
rect 603 15130 807 15140
rect 841 15130 1026 15164
rect 603 15106 1026 15130
rect 603 15072 632 15106
rect 666 15092 1026 15106
rect 666 15072 807 15092
rect 603 15058 807 15072
rect 841 15088 1026 15092
rect 13968 15195 14122 15229
rect 14156 15208 14297 15229
rect 14331 15208 14361 15242
rect 14156 15195 14361 15208
rect 13968 15174 14361 15195
rect 13968 15157 14297 15174
rect 13968 15123 14122 15157
rect 14156 15140 14297 15157
rect 14331 15140 14361 15174
rect 14156 15123 14361 15140
rect 13968 15106 14361 15123
rect 13968 15088 14297 15106
rect 841 15085 14297 15088
rect 841 15058 14122 15085
rect 603 15051 14122 15058
rect 14156 15072 14297 15085
rect 14331 15072 14361 15106
rect 14156 15051 14361 15072
rect 603 15038 14361 15051
rect 603 15004 632 15038
rect 666 15004 14297 15038
rect 14331 15004 14361 15038
rect 603 14970 14361 15004
rect 603 14936 632 14970
rect 666 14942 14297 14970
rect 666 14936 891 14942
rect 603 14908 891 14936
rect 925 14908 963 14942
rect 997 14908 1035 14942
rect 1069 14908 1107 14942
rect 1141 14908 1179 14942
rect 1213 14908 1251 14942
rect 1285 14908 1323 14942
rect 1357 14908 1395 14942
rect 1429 14908 1467 14942
rect 1501 14908 1539 14942
rect 1573 14908 1611 14942
rect 1645 14908 1683 14942
rect 1717 14908 1755 14942
rect 1789 14908 1827 14942
rect 1861 14908 1899 14942
rect 1933 14908 1971 14942
rect 2005 14908 2043 14942
rect 2077 14908 2115 14942
rect 2149 14908 2187 14942
rect 2221 14908 2259 14942
rect 2293 14908 2331 14942
rect 2365 14908 2403 14942
rect 2437 14908 2475 14942
rect 2509 14908 2547 14942
rect 2581 14908 2619 14942
rect 2653 14908 2691 14942
rect 2725 14908 2763 14942
rect 2797 14908 2835 14942
rect 2869 14908 2907 14942
rect 2941 14908 2979 14942
rect 3013 14908 3051 14942
rect 3085 14908 3123 14942
rect 3157 14908 3195 14942
rect 3229 14908 3267 14942
rect 3301 14908 3339 14942
rect 3373 14908 3411 14942
rect 3445 14908 3483 14942
rect 3517 14908 3555 14942
rect 3589 14908 3627 14942
rect 3661 14908 3699 14942
rect 3733 14908 3771 14942
rect 3805 14908 3843 14942
rect 3877 14908 3915 14942
rect 3949 14908 3987 14942
rect 4021 14908 4059 14942
rect 4093 14908 4131 14942
rect 4165 14908 4203 14942
rect 4237 14908 4275 14942
rect 4309 14908 4347 14942
rect 4381 14908 4419 14942
rect 4453 14908 4491 14942
rect 4525 14908 4563 14942
rect 4597 14908 4635 14942
rect 4669 14908 4707 14942
rect 4741 14908 4779 14942
rect 4813 14908 4851 14942
rect 4885 14908 4923 14942
rect 4957 14908 4995 14942
rect 5029 14908 5067 14942
rect 5101 14908 5139 14942
rect 5173 14908 5211 14942
rect 5245 14908 5283 14942
rect 5317 14908 5355 14942
rect 5389 14908 5427 14942
rect 5461 14908 5499 14942
rect 5533 14908 5571 14942
rect 5605 14908 5643 14942
rect 5677 14908 5715 14942
rect 5749 14908 5787 14942
rect 5821 14908 5859 14942
rect 5893 14908 5931 14942
rect 5965 14908 6003 14942
rect 6037 14908 6075 14942
rect 6109 14908 6147 14942
rect 6181 14908 6219 14942
rect 6253 14908 6291 14942
rect 6325 14908 6363 14942
rect 6397 14908 6435 14942
rect 6469 14908 6507 14942
rect 6541 14908 6579 14942
rect 6613 14908 6651 14942
rect 6685 14908 6723 14942
rect 6757 14908 6795 14942
rect 6829 14908 6867 14942
rect 6901 14908 6939 14942
rect 6973 14908 7011 14942
rect 7045 14908 7083 14942
rect 7117 14908 7155 14942
rect 7189 14908 7227 14942
rect 7261 14908 7299 14942
rect 7333 14908 7371 14942
rect 7405 14908 7443 14942
rect 7477 14908 7515 14942
rect 7549 14908 7587 14942
rect 7621 14908 7659 14942
rect 7693 14908 7731 14942
rect 7765 14908 7803 14942
rect 7837 14908 7875 14942
rect 7909 14908 7947 14942
rect 7981 14908 8019 14942
rect 8053 14908 8091 14942
rect 8125 14908 8163 14942
rect 8197 14908 8235 14942
rect 8269 14908 8307 14942
rect 8341 14908 8379 14942
rect 8413 14908 8451 14942
rect 8485 14908 8523 14942
rect 8557 14908 8595 14942
rect 8629 14908 8667 14942
rect 8701 14908 8739 14942
rect 8773 14908 8811 14942
rect 8845 14908 8883 14942
rect 8917 14908 8955 14942
rect 8989 14908 9027 14942
rect 9061 14908 9099 14942
rect 9133 14908 9171 14942
rect 9205 14908 9243 14942
rect 9277 14908 9315 14942
rect 9349 14908 9387 14942
rect 9421 14908 9459 14942
rect 9493 14908 9531 14942
rect 9565 14908 9603 14942
rect 9637 14908 9675 14942
rect 9709 14908 9747 14942
rect 9781 14908 9819 14942
rect 9853 14908 9891 14942
rect 9925 14908 9963 14942
rect 9997 14908 10035 14942
rect 10069 14908 10107 14942
rect 10141 14908 10179 14942
rect 10213 14908 10251 14942
rect 10285 14908 10323 14942
rect 10357 14908 10395 14942
rect 10429 14908 10467 14942
rect 10501 14908 10539 14942
rect 10573 14908 10611 14942
rect 10645 14908 10683 14942
rect 10717 14908 10755 14942
rect 10789 14908 10827 14942
rect 10861 14908 10899 14942
rect 10933 14908 10971 14942
rect 11005 14908 11043 14942
rect 11077 14908 11115 14942
rect 11149 14908 11187 14942
rect 11221 14908 11259 14942
rect 11293 14908 11331 14942
rect 11365 14908 11403 14942
rect 11437 14908 11475 14942
rect 11509 14908 11547 14942
rect 11581 14908 11619 14942
rect 11653 14908 11691 14942
rect 11725 14908 11763 14942
rect 11797 14908 11835 14942
rect 11869 14908 11907 14942
rect 11941 14908 11979 14942
rect 12013 14908 12051 14942
rect 12085 14908 12123 14942
rect 12157 14908 12195 14942
rect 12229 14908 12267 14942
rect 12301 14908 12339 14942
rect 12373 14908 12411 14942
rect 12445 14908 12483 14942
rect 12517 14908 12555 14942
rect 12589 14908 12627 14942
rect 12661 14908 12699 14942
rect 12733 14908 12771 14942
rect 12805 14908 12843 14942
rect 12877 14908 12915 14942
rect 12949 14908 12987 14942
rect 13021 14908 13059 14942
rect 13093 14908 13131 14942
rect 13165 14908 13203 14942
rect 13237 14908 13275 14942
rect 13309 14908 13347 14942
rect 13381 14908 13419 14942
rect 13453 14908 13491 14942
rect 13525 14908 13563 14942
rect 13597 14908 13635 14942
rect 13669 14908 13707 14942
rect 13741 14908 13779 14942
rect 13813 14908 13851 14942
rect 13885 14908 13923 14942
rect 13957 14908 13995 14942
rect 14029 14936 14297 14942
rect 14331 14936 14361 14970
rect 14029 14908 14361 14936
rect 603 14902 14361 14908
rect 603 14868 632 14902
rect 666 14868 14297 14902
rect 14331 14868 14361 14902
rect 603 14775 14361 14868
rect 603 14741 766 14775
rect 800 14741 834 14775
rect 868 14774 902 14775
rect 936 14774 970 14775
rect 1004 14774 1038 14775
rect 1072 14774 1106 14775
rect 1140 14774 1174 14775
rect 868 14741 883 14774
rect 936 14741 955 14774
rect 1004 14741 1027 14774
rect 1072 14741 1099 14774
rect 1140 14741 1171 14774
rect 1208 14741 1242 14775
rect 1276 14774 1310 14775
rect 1344 14774 1378 14775
rect 1412 14774 1446 14775
rect 1480 14774 1514 14775
rect 1548 14774 1582 14775
rect 1616 14774 1650 14775
rect 1684 14774 1718 14775
rect 1752 14774 1786 14775
rect 1820 14774 1854 14775
rect 1277 14741 1310 14774
rect 1349 14741 1378 14774
rect 1421 14741 1446 14774
rect 1493 14741 1514 14774
rect 1565 14741 1582 14774
rect 1637 14741 1650 14774
rect 1709 14741 1718 14774
rect 1781 14741 1786 14774
rect 1853 14741 1854 14774
rect 1888 14774 1922 14775
rect 1956 14774 1990 14775
rect 2024 14774 2058 14775
rect 1888 14741 1891 14774
rect 1956 14741 1963 14774
rect 2024 14741 2035 14774
rect 2092 14741 2126 14775
rect 2160 14741 2194 14775
rect 2228 14741 2262 14775
rect 2296 14741 2330 14775
rect 2364 14741 2398 14775
rect 2432 14741 2466 14775
rect 2500 14741 2534 14775
rect 2568 14741 2602 14775
rect 2636 14741 2670 14775
rect 2704 14741 2738 14775
rect 2772 14741 2806 14775
rect 2840 14741 2874 14775
rect 2908 14741 2942 14775
rect 2976 14741 3010 14775
rect 3044 14741 3078 14775
rect 3112 14741 3146 14775
rect 3180 14741 3214 14775
rect 3248 14741 3282 14775
rect 3316 14741 3350 14775
rect 3384 14741 3418 14775
rect 3452 14741 3486 14775
rect 3520 14741 3554 14775
rect 3588 14741 3622 14775
rect 3656 14741 3690 14775
rect 3724 14741 3758 14775
rect 3792 14741 3826 14775
rect 3860 14741 3894 14775
rect 3928 14741 3962 14775
rect 3996 14741 4030 14775
rect 4064 14741 4098 14775
rect 4132 14741 4166 14775
rect 4200 14741 4234 14775
rect 4268 14741 4302 14775
rect 4336 14741 4370 14775
rect 4404 14741 4438 14775
rect 4472 14741 4506 14775
rect 4540 14741 4574 14775
rect 4608 14741 4642 14775
rect 4676 14741 4710 14775
rect 4744 14741 4778 14775
rect 4812 14741 4846 14775
rect 4880 14741 4914 14775
rect 4948 14741 4982 14775
rect 5016 14741 5050 14775
rect 5084 14741 5118 14775
rect 5152 14741 5186 14775
rect 5220 14741 5254 14775
rect 5288 14741 5322 14775
rect 5356 14741 5390 14775
rect 5424 14741 5458 14775
rect 5492 14741 5526 14775
rect 5560 14741 5594 14775
rect 5628 14741 5662 14775
rect 5696 14741 5730 14775
rect 5764 14741 5798 14775
rect 5832 14741 5866 14775
rect 5900 14741 5934 14775
rect 5968 14741 6002 14775
rect 6036 14741 6070 14775
rect 6104 14741 6138 14775
rect 6172 14741 6206 14775
rect 6240 14741 6274 14775
rect 6308 14741 6342 14775
rect 6376 14741 6410 14775
rect 6444 14741 6478 14775
rect 6512 14741 6546 14775
rect 6580 14741 6614 14775
rect 6648 14741 6682 14775
rect 6716 14741 6750 14775
rect 6784 14741 6818 14775
rect 6852 14741 6886 14775
rect 6920 14741 6954 14775
rect 6988 14741 7022 14775
rect 7056 14741 7090 14775
rect 7124 14741 7158 14775
rect 7192 14741 7226 14775
rect 7260 14741 7294 14775
rect 7328 14741 7362 14775
rect 7396 14741 7430 14775
rect 7464 14741 7498 14775
rect 7532 14741 7566 14775
rect 7600 14741 7634 14775
rect 7668 14741 7702 14775
rect 7736 14741 7770 14775
rect 7804 14741 7838 14775
rect 7872 14741 7906 14775
rect 7940 14741 7974 14775
rect 8008 14741 8042 14775
rect 8076 14741 8110 14775
rect 8144 14741 8178 14775
rect 8212 14741 8246 14775
rect 8280 14741 8314 14775
rect 8348 14741 8382 14775
rect 8416 14741 8450 14775
rect 8484 14741 8518 14775
rect 8552 14741 8586 14775
rect 8620 14741 8654 14775
rect 8688 14741 8722 14775
rect 8756 14741 8790 14775
rect 8824 14741 8858 14775
rect 8892 14741 8926 14775
rect 8960 14741 8994 14775
rect 9028 14741 9062 14775
rect 9096 14741 9130 14775
rect 9164 14741 9198 14775
rect 9232 14741 9266 14775
rect 9300 14741 9334 14775
rect 9368 14741 9402 14775
rect 9436 14741 9470 14775
rect 9504 14741 9538 14775
rect 9572 14741 9606 14775
rect 9640 14741 9674 14775
rect 9708 14741 9742 14775
rect 9776 14741 9810 14775
rect 9844 14741 9878 14775
rect 9912 14741 9946 14775
rect 9980 14741 10014 14775
rect 10048 14741 10082 14775
rect 10116 14741 10150 14775
rect 10184 14741 10218 14775
rect 10252 14741 10286 14775
rect 10320 14741 10354 14775
rect 10388 14741 10422 14775
rect 10456 14741 10490 14775
rect 10524 14741 10558 14775
rect 10592 14741 10626 14775
rect 10660 14741 10694 14775
rect 10728 14741 10762 14775
rect 10796 14741 10830 14775
rect 10864 14741 10898 14775
rect 10932 14741 10966 14775
rect 11000 14741 11034 14775
rect 11068 14741 11102 14775
rect 11136 14741 11170 14775
rect 11204 14741 11238 14775
rect 11272 14741 11306 14775
rect 11340 14741 11374 14775
rect 11408 14741 11442 14775
rect 11476 14741 11510 14775
rect 11544 14741 11578 14775
rect 11612 14741 11646 14775
rect 11680 14741 11714 14775
rect 11748 14741 11782 14775
rect 11816 14741 11850 14775
rect 11884 14741 11918 14775
rect 11952 14741 11986 14775
rect 12020 14741 12054 14775
rect 12088 14741 12122 14775
rect 12156 14741 12190 14775
rect 12224 14741 12258 14775
rect 12292 14741 12326 14775
rect 12360 14741 12394 14775
rect 12428 14741 12462 14775
rect 12496 14741 12530 14775
rect 12564 14741 12598 14775
rect 12632 14741 12666 14775
rect 12700 14741 12734 14775
rect 12768 14741 12802 14775
rect 12836 14741 12870 14775
rect 12904 14774 12938 14775
rect 12972 14774 13006 14775
rect 13040 14774 13074 14775
rect 13108 14774 13142 14775
rect 13176 14774 13210 14775
rect 13244 14774 13278 14775
rect 12917 14741 12938 14774
rect 12989 14741 13006 14774
rect 13061 14741 13074 14774
rect 13133 14741 13142 14774
rect 13205 14741 13210 14774
rect 13277 14741 13278 14774
rect 13312 14774 13346 14775
rect 13380 14774 13414 14775
rect 13448 14774 13482 14775
rect 13516 14774 13550 14775
rect 13584 14774 13618 14775
rect 13652 14774 13686 14775
rect 13720 14774 13754 14775
rect 13788 14774 13822 14775
rect 13312 14741 13315 14774
rect 13380 14741 13387 14774
rect 13448 14741 13459 14774
rect 13516 14741 13531 14774
rect 13584 14741 13603 14774
rect 13652 14741 13675 14774
rect 13720 14741 13747 14774
rect 13788 14741 13819 14774
rect 13856 14741 13890 14775
rect 13924 14774 13958 14775
rect 13992 14774 14026 14775
rect 14060 14774 14094 14775
rect 13925 14741 13958 14774
rect 13997 14741 14026 14774
rect 14069 14741 14094 14774
rect 14128 14741 14162 14775
rect 14196 14741 14361 14775
rect 603 14740 883 14741
rect 917 14740 955 14741
rect 989 14740 1027 14741
rect 1061 14740 1099 14741
rect 1133 14740 1171 14741
rect 1205 14740 1243 14741
rect 1277 14740 1315 14741
rect 1349 14740 1387 14741
rect 1421 14740 1459 14741
rect 1493 14740 1531 14741
rect 1565 14740 1603 14741
rect 1637 14740 1675 14741
rect 1709 14740 1747 14741
rect 1781 14740 1819 14741
rect 1853 14740 1891 14741
rect 1925 14740 1963 14741
rect 1997 14740 2035 14741
rect 2069 14740 12883 14741
rect 12917 14740 12955 14741
rect 12989 14740 13027 14741
rect 13061 14740 13099 14741
rect 13133 14740 13171 14741
rect 13205 14740 13243 14741
rect 13277 14740 13315 14741
rect 13349 14740 13387 14741
rect 13421 14740 13459 14741
rect 13493 14740 13531 14741
rect 13565 14740 13603 14741
rect 13637 14740 13675 14741
rect 13709 14740 13747 14741
rect 13781 14740 13819 14741
rect 13853 14740 13891 14741
rect 13925 14740 13963 14741
rect 13997 14740 14035 14741
rect 14069 14740 14361 14741
rect 603 14711 14361 14740
rect 14539 36192 14607 36226
rect 14641 36206 14724 36226
rect 14539 36172 14614 36192
rect 14648 36172 14724 36206
rect 14539 36158 14724 36172
rect 14539 36124 14607 36158
rect 14641 36134 14724 36158
rect 14539 36100 14614 36124
rect 14648 36100 14724 36134
rect 14539 36090 14724 36100
rect 14539 36056 14607 36090
rect 14641 36062 14724 36090
rect 14539 36028 14614 36056
rect 14648 36028 14724 36062
rect 14539 36022 14724 36028
rect 14539 35988 14607 36022
rect 14641 35990 14724 36022
rect 14539 35956 14614 35988
rect 14648 35956 14724 35990
rect 14539 35954 14724 35956
rect 14539 35920 14607 35954
rect 14641 35920 14724 35954
rect 14539 35918 14724 35920
rect 14539 35886 14614 35918
rect 14539 35852 14607 35886
rect 14648 35884 14724 35918
rect 14641 35852 14724 35884
rect 14539 35846 14724 35852
rect 14539 35818 14614 35846
rect 14539 35784 14607 35818
rect 14648 35812 14724 35846
rect 14641 35784 14724 35812
rect 14539 35774 14724 35784
rect 14539 35750 14614 35774
rect 14539 35716 14607 35750
rect 14648 35740 14724 35774
rect 14641 35716 14724 35740
rect 14539 35702 14724 35716
rect 14539 35682 14614 35702
rect 14539 35648 14607 35682
rect 14648 35668 14724 35702
rect 14641 35648 14724 35668
rect 14539 35630 14724 35648
rect 14539 35614 14614 35630
rect 14539 35580 14607 35614
rect 14648 35596 14724 35630
rect 14641 35580 14724 35596
rect 14539 35558 14724 35580
rect 14539 35546 14614 35558
rect 14539 35512 14607 35546
rect 14648 35524 14724 35558
rect 14641 35512 14724 35524
rect 14539 35486 14724 35512
rect 14539 35478 14614 35486
rect 14539 35444 14607 35478
rect 14648 35452 14724 35486
rect 14641 35444 14724 35452
rect 14539 35414 14724 35444
rect 14539 35410 14614 35414
rect 14539 35376 14607 35410
rect 14648 35380 14724 35414
rect 14641 35376 14724 35380
rect 14539 35342 14724 35376
rect 14539 35308 14607 35342
rect 14648 35308 14724 35342
rect 14539 35274 14724 35308
rect 14539 35240 14607 35274
rect 14641 35270 14724 35274
rect 14539 35236 14614 35240
rect 14648 35236 14724 35270
rect 14539 35206 14724 35236
rect 14539 35172 14607 35206
rect 14641 35198 14724 35206
rect 14539 35164 14614 35172
rect 14648 35164 14724 35198
rect 14539 35138 14724 35164
rect 14539 35104 14607 35138
rect 14641 35126 14724 35138
rect 14539 35092 14614 35104
rect 14648 35092 14724 35126
rect 14539 35070 14724 35092
rect 14539 35036 14607 35070
rect 14641 35054 14724 35070
rect 14539 35020 14614 35036
rect 14648 35020 14724 35054
rect 14539 35002 14724 35020
rect 14539 34968 14607 35002
rect 14641 34982 14724 35002
rect 14539 34948 14614 34968
rect 14648 34948 14724 34982
rect 14539 34934 14724 34948
rect 14539 34900 14607 34934
rect 14641 34910 14724 34934
rect 14539 34876 14614 34900
rect 14648 34876 14724 34910
rect 14539 34866 14724 34876
rect 14539 34832 14607 34866
rect 14641 34838 14724 34866
rect 14539 34804 14614 34832
rect 14648 34804 14724 34838
rect 14539 34798 14724 34804
rect 14539 34764 14607 34798
rect 14641 34766 14724 34798
rect 14539 34732 14614 34764
rect 14648 34732 14724 34766
rect 14539 34730 14724 34732
rect 14539 34696 14607 34730
rect 14641 34696 14724 34730
rect 14539 34694 14724 34696
rect 14539 34662 14614 34694
rect 14539 34628 14607 34662
rect 14648 34660 14724 34694
rect 14641 34628 14724 34660
rect 14539 34622 14724 34628
rect 14539 34594 14614 34622
rect 14539 34560 14607 34594
rect 14648 34588 14724 34622
rect 14641 34560 14724 34588
rect 14539 34550 14724 34560
rect 14539 34526 14614 34550
rect 14539 34492 14607 34526
rect 14648 34516 14724 34550
rect 14641 34492 14724 34516
rect 14539 34478 14724 34492
rect 14539 34458 14614 34478
rect 14539 34424 14607 34458
rect 14648 34444 14724 34478
rect 14641 34424 14724 34444
rect 14539 34406 14724 34424
rect 14539 34390 14614 34406
rect 14539 34356 14607 34390
rect 14648 34372 14724 34406
rect 14641 34356 14724 34372
rect 14539 34334 14724 34356
rect 14539 34322 14614 34334
rect 14539 34288 14607 34322
rect 14648 34300 14724 34334
rect 14641 34288 14724 34300
rect 14539 34262 14724 34288
rect 14539 34254 14614 34262
rect 14539 34220 14607 34254
rect 14648 34228 14724 34262
rect 14641 34220 14724 34228
rect 14539 34190 14724 34220
rect 14539 34186 14614 34190
rect 14539 34152 14607 34186
rect 14648 34156 14724 34190
rect 14641 34152 14724 34156
rect 14539 34118 14724 34152
rect 14539 34084 14607 34118
rect 14648 34084 14724 34118
rect 14539 34050 14724 34084
rect 14539 34016 14607 34050
rect 14641 34046 14724 34050
rect 14539 34012 14614 34016
rect 14648 34012 14724 34046
rect 14539 33982 14724 34012
rect 14539 33948 14607 33982
rect 14641 33974 14724 33982
rect 14539 33940 14614 33948
rect 14648 33940 14724 33974
rect 14539 33914 14724 33940
rect 14539 33880 14607 33914
rect 14641 33902 14724 33914
rect 14539 33868 14614 33880
rect 14648 33868 14724 33902
rect 14539 33846 14724 33868
rect 14539 33812 14607 33846
rect 14641 33830 14724 33846
rect 14539 33796 14614 33812
rect 14648 33796 14724 33830
rect 14539 33778 14724 33796
rect 14539 33744 14607 33778
rect 14641 33758 14724 33778
rect 14539 33724 14614 33744
rect 14648 33724 14724 33758
rect 14539 33710 14724 33724
rect 14539 33676 14607 33710
rect 14641 33686 14724 33710
rect 14539 33652 14614 33676
rect 14648 33652 14724 33686
rect 14539 33642 14724 33652
rect 14539 33608 14607 33642
rect 14641 33614 14724 33642
rect 14539 33580 14614 33608
rect 14648 33580 14724 33614
rect 14539 33574 14724 33580
rect 14539 33540 14607 33574
rect 14641 33542 14724 33574
rect 14539 33508 14614 33540
rect 14648 33508 14724 33542
rect 14539 33506 14724 33508
rect 14539 33472 14607 33506
rect 14641 33472 14724 33506
rect 14539 33470 14724 33472
rect 14539 33438 14614 33470
rect 14539 33404 14607 33438
rect 14648 33436 14724 33470
rect 14641 33404 14724 33436
rect 14539 33398 14724 33404
rect 14539 33370 14614 33398
rect 14539 33336 14607 33370
rect 14648 33364 14724 33398
rect 14641 33336 14724 33364
rect 14539 33326 14724 33336
rect 14539 33302 14614 33326
rect 14539 33268 14607 33302
rect 14648 33292 14724 33326
rect 14641 33268 14724 33292
rect 14539 33254 14724 33268
rect 14539 33234 14614 33254
rect 14539 33200 14607 33234
rect 14648 33220 14724 33254
rect 14641 33200 14724 33220
rect 14539 33182 14724 33200
rect 14539 33166 14614 33182
rect 14539 33132 14607 33166
rect 14648 33148 14724 33182
rect 14641 33132 14724 33148
rect 14539 33110 14724 33132
rect 14539 33098 14614 33110
rect 14539 33064 14607 33098
rect 14648 33076 14724 33110
rect 14641 33064 14724 33076
rect 14539 33038 14724 33064
rect 14539 33030 14614 33038
rect 14539 32996 14607 33030
rect 14648 33004 14724 33038
rect 14641 32996 14724 33004
rect 14539 32966 14724 32996
rect 14539 32962 14614 32966
rect 14539 32928 14607 32962
rect 14648 32932 14724 32966
rect 14641 32928 14724 32932
rect 14539 32894 14724 32928
rect 14539 32860 14607 32894
rect 14648 32860 14724 32894
rect 14539 32826 14724 32860
rect 14539 32792 14607 32826
rect 14641 32822 14724 32826
rect 14539 32788 14614 32792
rect 14648 32788 14724 32822
rect 14539 32758 14724 32788
rect 14539 32724 14607 32758
rect 14641 32750 14724 32758
rect 14539 32716 14614 32724
rect 14648 32716 14724 32750
rect 14539 32690 14724 32716
rect 14539 32656 14607 32690
rect 14641 32678 14724 32690
rect 14539 32644 14614 32656
rect 14648 32644 14724 32678
rect 14539 32622 14724 32644
rect 14539 32588 14607 32622
rect 14641 32606 14724 32622
rect 14539 32572 14614 32588
rect 14648 32572 14724 32606
rect 14539 32554 14724 32572
rect 14539 32520 14607 32554
rect 14641 32534 14724 32554
rect 14539 32500 14614 32520
rect 14648 32500 14724 32534
rect 14539 32486 14724 32500
rect 14539 32452 14607 32486
rect 14641 32462 14724 32486
rect 14539 32428 14614 32452
rect 14648 32428 14724 32462
rect 14539 32418 14724 32428
rect 14539 32384 14607 32418
rect 14641 32390 14724 32418
rect 14539 32356 14614 32384
rect 14648 32356 14724 32390
rect 14539 32350 14724 32356
rect 14539 32316 14607 32350
rect 14641 32318 14724 32350
rect 14539 32284 14614 32316
rect 14648 32284 14724 32318
rect 14539 32282 14724 32284
rect 14539 32248 14607 32282
rect 14641 32248 14724 32282
rect 14539 32246 14724 32248
rect 14539 32214 14614 32246
rect 14539 32180 14607 32214
rect 14648 32212 14724 32246
rect 14641 32180 14724 32212
rect 14539 32174 14724 32180
rect 14539 32146 14614 32174
rect 14539 32112 14607 32146
rect 14648 32140 14724 32174
rect 14641 32112 14724 32140
rect 14539 32102 14724 32112
rect 14539 32078 14614 32102
rect 14539 32044 14607 32078
rect 14648 32068 14724 32102
rect 14641 32044 14724 32068
rect 14539 32030 14724 32044
rect 14539 32010 14614 32030
rect 14539 31976 14607 32010
rect 14648 31996 14724 32030
rect 14641 31976 14724 31996
rect 14539 31958 14724 31976
rect 14539 31942 14614 31958
rect 14539 31908 14607 31942
rect 14648 31924 14724 31958
rect 14641 31908 14724 31924
rect 14539 31886 14724 31908
rect 14539 31874 14614 31886
rect 14539 31840 14607 31874
rect 14648 31852 14724 31886
rect 14641 31840 14724 31852
rect 14539 31814 14724 31840
rect 14539 31806 14614 31814
rect 14539 31772 14607 31806
rect 14648 31780 14724 31814
rect 14641 31772 14724 31780
rect 14539 31742 14724 31772
rect 14539 31738 14614 31742
rect 14539 31704 14607 31738
rect 14648 31708 14724 31742
rect 14641 31704 14724 31708
rect 14539 31670 14724 31704
rect 14539 31636 14607 31670
rect 14648 31636 14724 31670
rect 14539 31602 14724 31636
rect 14539 31568 14607 31602
rect 14641 31598 14724 31602
rect 14539 31564 14614 31568
rect 14648 31564 14724 31598
rect 14539 31534 14724 31564
rect 14539 31500 14607 31534
rect 14641 31526 14724 31534
rect 14539 31492 14614 31500
rect 14648 31492 14724 31526
rect 14539 31466 14724 31492
rect 14539 31432 14607 31466
rect 14641 31454 14724 31466
rect 14539 31420 14614 31432
rect 14648 31420 14724 31454
rect 14539 31398 14724 31420
rect 14539 31364 14607 31398
rect 14641 31382 14724 31398
rect 14539 31348 14614 31364
rect 14648 31348 14724 31382
rect 14539 31330 14724 31348
rect 14539 31296 14607 31330
rect 14641 31310 14724 31330
rect 14539 31276 14614 31296
rect 14648 31276 14724 31310
rect 14539 31262 14724 31276
rect 14539 31228 14607 31262
rect 14641 31238 14724 31262
rect 14539 31204 14614 31228
rect 14648 31204 14724 31238
rect 14539 31194 14724 31204
rect 14539 31160 14607 31194
rect 14641 31166 14724 31194
rect 14539 31132 14614 31160
rect 14648 31132 14724 31166
rect 14539 31126 14724 31132
rect 14539 31092 14607 31126
rect 14641 31094 14724 31126
rect 14539 31060 14614 31092
rect 14648 31060 14724 31094
rect 14539 31058 14724 31060
rect 14539 31024 14607 31058
rect 14641 31024 14724 31058
rect 14539 31022 14724 31024
rect 14539 30990 14614 31022
rect 14539 30956 14607 30990
rect 14648 30988 14724 31022
rect 14641 30956 14724 30988
rect 14539 30950 14724 30956
rect 14539 30922 14614 30950
rect 14539 30888 14607 30922
rect 14648 30916 14724 30950
rect 14641 30888 14724 30916
rect 14539 30878 14724 30888
rect 14539 30854 14614 30878
rect 14539 30820 14607 30854
rect 14648 30844 14724 30878
rect 14641 30820 14724 30844
rect 14539 30806 14724 30820
rect 14539 30786 14614 30806
rect 14539 30752 14607 30786
rect 14648 30772 14724 30806
rect 14641 30752 14724 30772
rect 14539 30734 14724 30752
rect 14539 30718 14614 30734
rect 14539 30684 14607 30718
rect 14648 30700 14724 30734
rect 14641 30684 14724 30700
rect 14539 30662 14724 30684
rect 14539 30650 14614 30662
rect 14539 30616 14607 30650
rect 14648 30628 14724 30662
rect 14641 30616 14724 30628
rect 14539 30590 14724 30616
rect 14539 30582 14614 30590
rect 14539 30548 14607 30582
rect 14648 30556 14724 30590
rect 14641 30548 14724 30556
rect 14539 30518 14724 30548
rect 14539 30514 14614 30518
rect 14539 30480 14607 30514
rect 14648 30484 14724 30518
rect 14641 30480 14724 30484
rect 14539 30446 14724 30480
rect 14539 30412 14607 30446
rect 14648 30412 14724 30446
rect 14539 30378 14724 30412
rect 14539 30344 14607 30378
rect 14641 30374 14724 30378
rect 14539 30340 14614 30344
rect 14648 30340 14724 30374
rect 14539 30310 14724 30340
rect 14539 30276 14607 30310
rect 14641 30302 14724 30310
rect 14539 30268 14614 30276
rect 14648 30268 14724 30302
rect 14539 30242 14724 30268
rect 14539 30208 14607 30242
rect 14641 30230 14724 30242
rect 14539 30196 14614 30208
rect 14648 30196 14724 30230
rect 14539 30174 14724 30196
rect 14539 30140 14607 30174
rect 14641 30158 14724 30174
rect 14539 30124 14614 30140
rect 14648 30124 14724 30158
rect 14539 30106 14724 30124
rect 14539 30072 14607 30106
rect 14641 30086 14724 30106
rect 14539 30052 14614 30072
rect 14648 30052 14724 30086
rect 14539 30038 14724 30052
rect 14539 30004 14607 30038
rect 14641 30014 14724 30038
rect 14539 29980 14614 30004
rect 14648 29980 14724 30014
rect 14539 29970 14724 29980
rect 14539 29936 14607 29970
rect 14641 29942 14724 29970
rect 14539 29908 14614 29936
rect 14648 29908 14724 29942
rect 14539 29902 14724 29908
rect 14539 29868 14607 29902
rect 14641 29870 14724 29902
rect 14539 29836 14614 29868
rect 14648 29836 14724 29870
rect 14539 29834 14724 29836
rect 14539 29800 14607 29834
rect 14641 29800 14724 29834
rect 14539 29798 14724 29800
rect 14539 29766 14614 29798
rect 14539 29732 14607 29766
rect 14648 29764 14724 29798
rect 14641 29732 14724 29764
rect 14539 29726 14724 29732
rect 14539 29698 14614 29726
rect 14539 29664 14607 29698
rect 14648 29692 14724 29726
rect 14641 29664 14724 29692
rect 14539 29654 14724 29664
rect 14539 29630 14614 29654
rect 14539 29596 14607 29630
rect 14648 29620 14724 29654
rect 14641 29596 14724 29620
rect 14539 29582 14724 29596
rect 14539 29562 14614 29582
rect 14539 29528 14607 29562
rect 14648 29548 14724 29582
rect 14641 29528 14724 29548
rect 14539 29510 14724 29528
rect 14539 29494 14614 29510
rect 14539 29460 14607 29494
rect 14648 29476 14724 29510
rect 14641 29460 14724 29476
rect 14539 29438 14724 29460
rect 14539 29426 14614 29438
rect 14539 29392 14607 29426
rect 14648 29404 14724 29438
rect 14641 29392 14724 29404
rect 14539 29366 14724 29392
rect 14539 29358 14614 29366
rect 14539 29324 14607 29358
rect 14648 29332 14724 29366
rect 14641 29324 14724 29332
rect 14539 29294 14724 29324
rect 14539 29290 14614 29294
rect 14539 29256 14607 29290
rect 14648 29260 14724 29294
rect 14641 29256 14724 29260
rect 14539 29222 14724 29256
rect 14539 29188 14607 29222
rect 14648 29188 14724 29222
rect 14539 29154 14724 29188
rect 14539 29120 14607 29154
rect 14641 29150 14724 29154
rect 14539 29116 14614 29120
rect 14648 29116 14724 29150
rect 14539 29086 14724 29116
rect 14539 29052 14607 29086
rect 14641 29078 14724 29086
rect 14539 29044 14614 29052
rect 14648 29044 14724 29078
rect 14539 29018 14724 29044
rect 14539 28984 14607 29018
rect 14641 29006 14724 29018
rect 14539 28972 14614 28984
rect 14648 28972 14724 29006
rect 14539 28950 14724 28972
rect 14539 28916 14607 28950
rect 14641 28934 14724 28950
rect 14539 28900 14614 28916
rect 14648 28900 14724 28934
rect 14539 28882 14724 28900
rect 14539 28848 14607 28882
rect 14641 28862 14724 28882
rect 14539 28828 14614 28848
rect 14648 28828 14724 28862
rect 14539 28814 14724 28828
rect 14539 28780 14607 28814
rect 14641 28790 14724 28814
rect 14539 28756 14614 28780
rect 14648 28756 14724 28790
rect 14539 28746 14724 28756
rect 14539 28712 14607 28746
rect 14641 28718 14724 28746
rect 14539 28684 14614 28712
rect 14648 28684 14724 28718
rect 14539 28678 14724 28684
rect 14539 28644 14607 28678
rect 14641 28646 14724 28678
rect 14539 28612 14614 28644
rect 14648 28612 14724 28646
rect 14539 28610 14724 28612
rect 14539 28576 14607 28610
rect 14641 28576 14724 28610
rect 14539 28574 14724 28576
rect 14539 28542 14614 28574
rect 14539 28508 14607 28542
rect 14648 28540 14724 28574
rect 14641 28508 14724 28540
rect 14539 28502 14724 28508
rect 14539 28474 14614 28502
rect 14539 28440 14607 28474
rect 14648 28468 14724 28502
rect 14641 28440 14724 28468
rect 14539 28430 14724 28440
rect 14539 28406 14614 28430
rect 14539 28372 14607 28406
rect 14648 28396 14724 28430
rect 14641 28372 14724 28396
rect 14539 28358 14724 28372
rect 14539 28338 14614 28358
rect 14539 28304 14607 28338
rect 14648 28324 14724 28358
rect 14641 28304 14724 28324
rect 14539 28286 14724 28304
rect 14539 28270 14614 28286
rect 14539 28236 14607 28270
rect 14648 28252 14724 28286
rect 14641 28236 14724 28252
rect 14539 28214 14724 28236
rect 14539 28202 14614 28214
rect 14539 28168 14607 28202
rect 14648 28180 14724 28214
rect 14641 28168 14724 28180
rect 14539 28142 14724 28168
rect 14539 28134 14614 28142
rect 14539 28100 14607 28134
rect 14648 28108 14724 28142
rect 14641 28100 14724 28108
rect 14539 28070 14724 28100
rect 14539 28066 14614 28070
rect 14539 28032 14607 28066
rect 14648 28036 14724 28070
rect 14641 28032 14724 28036
rect 14539 27998 14724 28032
rect 14539 27964 14607 27998
rect 14648 27964 14724 27998
rect 14539 27930 14724 27964
rect 14539 27896 14607 27930
rect 14641 27926 14724 27930
rect 14539 27892 14614 27896
rect 14648 27892 14724 27926
rect 14539 27862 14724 27892
rect 14539 27828 14607 27862
rect 14641 27854 14724 27862
rect 14539 27820 14614 27828
rect 14648 27820 14724 27854
rect 14539 27794 14724 27820
rect 14539 27760 14607 27794
rect 14641 27782 14724 27794
rect 14539 27748 14614 27760
rect 14648 27748 14724 27782
rect 14539 27726 14724 27748
rect 14539 27692 14607 27726
rect 14641 27710 14724 27726
rect 14539 27676 14614 27692
rect 14648 27676 14724 27710
rect 14539 27658 14724 27676
rect 14539 27624 14607 27658
rect 14641 27638 14724 27658
rect 14539 27604 14614 27624
rect 14648 27604 14724 27638
rect 14539 27590 14724 27604
rect 14539 27556 14607 27590
rect 14641 27566 14724 27590
rect 14539 27532 14614 27556
rect 14648 27532 14724 27566
rect 14539 27522 14724 27532
rect 14539 27488 14607 27522
rect 14641 27494 14724 27522
rect 14539 27460 14614 27488
rect 14648 27460 14724 27494
rect 14539 27454 14724 27460
rect 14539 27420 14607 27454
rect 14641 27422 14724 27454
rect 14539 27388 14614 27420
rect 14648 27388 14724 27422
rect 14539 27386 14724 27388
rect 14539 27352 14607 27386
rect 14641 27352 14724 27386
rect 14539 27350 14724 27352
rect 14539 27318 14614 27350
rect 14539 27284 14607 27318
rect 14648 27316 14724 27350
rect 14641 27284 14724 27316
rect 14539 27278 14724 27284
rect 14539 27250 14614 27278
rect 14539 27216 14607 27250
rect 14648 27244 14724 27278
rect 14641 27216 14724 27244
rect 14539 27206 14724 27216
rect 14539 27182 14614 27206
rect 14539 27148 14607 27182
rect 14648 27172 14724 27206
rect 14641 27148 14724 27172
rect 14539 27134 14724 27148
rect 14539 27114 14614 27134
rect 14539 27080 14607 27114
rect 14648 27100 14724 27134
rect 14641 27080 14724 27100
rect 14539 27062 14724 27080
rect 14539 27046 14614 27062
rect 14539 27012 14607 27046
rect 14648 27028 14724 27062
rect 14641 27012 14724 27028
rect 14539 26990 14724 27012
rect 14539 26978 14614 26990
rect 14539 26944 14607 26978
rect 14648 26956 14724 26990
rect 14641 26944 14724 26956
rect 14539 26918 14724 26944
rect 14539 26910 14614 26918
rect 14539 26876 14607 26910
rect 14648 26884 14724 26918
rect 14641 26876 14724 26884
rect 14539 26846 14724 26876
rect 14539 26842 14614 26846
rect 14539 26808 14607 26842
rect 14648 26812 14724 26846
rect 14641 26808 14724 26812
rect 14539 26774 14724 26808
rect 14539 26740 14607 26774
rect 14648 26740 14724 26774
rect 14539 26706 14724 26740
rect 14539 26672 14607 26706
rect 14641 26702 14724 26706
rect 14539 26668 14614 26672
rect 14648 26668 14724 26702
rect 14539 26638 14724 26668
rect 14539 26604 14607 26638
rect 14641 26630 14724 26638
rect 14539 26596 14614 26604
rect 14648 26596 14724 26630
rect 14539 26570 14724 26596
rect 14539 26536 14607 26570
rect 14641 26558 14724 26570
rect 14539 26524 14614 26536
rect 14648 26524 14724 26558
rect 14539 26502 14724 26524
rect 14539 26468 14607 26502
rect 14641 26486 14724 26502
rect 14539 26452 14614 26468
rect 14648 26452 14724 26486
rect 14539 26434 14724 26452
rect 14539 26400 14607 26434
rect 14641 26414 14724 26434
rect 14539 26380 14614 26400
rect 14648 26380 14724 26414
rect 14539 26366 14724 26380
rect 14539 26332 14607 26366
rect 14641 26342 14724 26366
rect 14539 26308 14614 26332
rect 14648 26308 14724 26342
rect 14539 26298 14724 26308
rect 14539 26264 14607 26298
rect 14641 26270 14724 26298
rect 14539 26236 14614 26264
rect 14648 26236 14724 26270
rect 14539 26230 14724 26236
rect 14539 26196 14607 26230
rect 14641 26198 14724 26230
rect 14539 26164 14614 26196
rect 14648 26164 14724 26198
rect 14539 26162 14724 26164
rect 14539 26128 14607 26162
rect 14641 26128 14724 26162
rect 14539 26126 14724 26128
rect 14539 26094 14614 26126
rect 14539 26060 14607 26094
rect 14648 26092 14724 26126
rect 14641 26060 14724 26092
rect 14539 26054 14724 26060
rect 14539 26026 14614 26054
rect 14539 25992 14607 26026
rect 14648 26020 14724 26054
rect 14641 25992 14724 26020
rect 14539 25982 14724 25992
rect 14539 25958 14614 25982
rect 14539 25924 14607 25958
rect 14648 25948 14724 25982
rect 14641 25924 14724 25948
rect 14539 25910 14724 25924
rect 14539 25890 14614 25910
rect 14539 25856 14607 25890
rect 14648 25876 14724 25910
rect 14641 25856 14724 25876
rect 14539 25838 14724 25856
rect 14539 25822 14614 25838
rect 14539 25788 14607 25822
rect 14648 25804 14724 25838
rect 14641 25788 14724 25804
rect 14539 25766 14724 25788
rect 14539 25754 14614 25766
rect 14539 25720 14607 25754
rect 14648 25732 14724 25766
rect 14641 25720 14724 25732
rect 14539 25694 14724 25720
rect 14539 25686 14614 25694
rect 14539 25652 14607 25686
rect 14648 25660 14724 25694
rect 14641 25652 14724 25660
rect 14539 25622 14724 25652
rect 14539 25618 14614 25622
rect 14539 25584 14607 25618
rect 14648 25588 14724 25622
rect 14641 25584 14724 25588
rect 14539 25550 14724 25584
rect 14539 25516 14607 25550
rect 14648 25516 14724 25550
rect 14539 25482 14724 25516
rect 14539 25448 14607 25482
rect 14641 25478 14724 25482
rect 14539 25444 14614 25448
rect 14648 25444 14724 25478
rect 14539 25414 14724 25444
rect 14539 25380 14607 25414
rect 14641 25406 14724 25414
rect 14539 25372 14614 25380
rect 14648 25372 14724 25406
rect 14539 25346 14724 25372
rect 14539 25312 14607 25346
rect 14641 25334 14724 25346
rect 14539 25300 14614 25312
rect 14648 25300 14724 25334
rect 14539 25278 14724 25300
rect 14539 25244 14607 25278
rect 14641 25262 14724 25278
rect 14539 25228 14614 25244
rect 14648 25228 14724 25262
rect 14539 25210 14724 25228
rect 14539 25176 14607 25210
rect 14641 25190 14724 25210
rect 14539 25156 14614 25176
rect 14648 25156 14724 25190
rect 14539 25142 14724 25156
rect 14539 25108 14607 25142
rect 14641 25118 14724 25142
rect 14539 25084 14614 25108
rect 14648 25084 14724 25118
rect 14539 25074 14724 25084
rect 14539 25040 14607 25074
rect 14641 25046 14724 25074
rect 14539 25012 14614 25040
rect 14648 25012 14724 25046
rect 14539 25006 14724 25012
rect 14539 24972 14607 25006
rect 14641 24974 14724 25006
rect 14539 24940 14614 24972
rect 14648 24940 14724 24974
rect 14539 24938 14724 24940
rect 14539 24904 14607 24938
rect 14641 24904 14724 24938
rect 14539 24902 14724 24904
rect 14539 24870 14614 24902
rect 14539 24836 14607 24870
rect 14648 24868 14724 24902
rect 14641 24836 14724 24868
rect 14539 24830 14724 24836
rect 14539 24802 14614 24830
rect 14539 24768 14607 24802
rect 14648 24796 14724 24830
rect 14641 24768 14724 24796
rect 14539 24758 14724 24768
rect 14539 24734 14614 24758
rect 14539 24700 14607 24734
rect 14648 24724 14724 24758
rect 14641 24700 14724 24724
rect 14539 24686 14724 24700
rect 14539 24666 14614 24686
rect 14539 24632 14607 24666
rect 14648 24652 14724 24686
rect 14641 24632 14724 24652
rect 14539 24614 14724 24632
rect 14539 24598 14614 24614
rect 14539 24564 14607 24598
rect 14648 24580 14724 24614
rect 14641 24564 14724 24580
rect 14539 24542 14724 24564
rect 14539 24530 14614 24542
rect 14539 24496 14607 24530
rect 14648 24508 14724 24542
rect 14641 24496 14724 24508
rect 14539 24470 14724 24496
rect 14539 24462 14614 24470
rect 14539 24428 14607 24462
rect 14648 24436 14724 24470
rect 14641 24428 14724 24436
rect 14539 24398 14724 24428
rect 14539 24394 14614 24398
rect 14539 24360 14607 24394
rect 14648 24364 14724 24398
rect 14641 24360 14724 24364
rect 14539 24326 14724 24360
rect 14539 24292 14607 24326
rect 14648 24292 14724 24326
rect 14539 24258 14724 24292
rect 14539 24224 14607 24258
rect 14641 24254 14724 24258
rect 14539 24220 14614 24224
rect 14648 24220 14724 24254
rect 14539 24190 14724 24220
rect 14539 24156 14607 24190
rect 14641 24182 14724 24190
rect 14539 24148 14614 24156
rect 14648 24148 14724 24182
rect 14539 24122 14724 24148
rect 14539 24088 14607 24122
rect 14641 24110 14724 24122
rect 14539 24076 14614 24088
rect 14648 24076 14724 24110
rect 14539 24054 14724 24076
rect 14539 24020 14607 24054
rect 14641 24038 14724 24054
rect 14539 24004 14614 24020
rect 14648 24004 14724 24038
rect 14539 23986 14724 24004
rect 14539 23952 14607 23986
rect 14641 23966 14724 23986
rect 14539 23932 14614 23952
rect 14648 23932 14724 23966
rect 14539 23918 14724 23932
rect 14539 23884 14607 23918
rect 14641 23894 14724 23918
rect 14539 23860 14614 23884
rect 14648 23860 14724 23894
rect 14539 23850 14724 23860
rect 14539 23816 14607 23850
rect 14641 23822 14724 23850
rect 14539 23788 14614 23816
rect 14648 23788 14724 23822
rect 14539 23782 14724 23788
rect 14539 23748 14607 23782
rect 14641 23750 14724 23782
rect 14539 23716 14614 23748
rect 14648 23716 14724 23750
rect 14539 23714 14724 23716
rect 14539 23680 14607 23714
rect 14641 23680 14724 23714
rect 14539 23678 14724 23680
rect 14539 23646 14614 23678
rect 14539 23612 14607 23646
rect 14648 23644 14724 23678
rect 14641 23612 14724 23644
rect 14539 23606 14724 23612
rect 14539 23578 14614 23606
rect 14539 23544 14607 23578
rect 14648 23572 14724 23606
rect 14641 23544 14724 23572
rect 14539 23534 14724 23544
rect 14539 23510 14614 23534
rect 14539 23476 14607 23510
rect 14648 23500 14724 23534
rect 14641 23476 14724 23500
rect 14539 23462 14724 23476
rect 14539 23442 14614 23462
rect 14539 23408 14607 23442
rect 14648 23428 14724 23462
rect 14641 23408 14724 23428
rect 14539 23390 14724 23408
rect 14539 23374 14614 23390
rect 14539 23340 14607 23374
rect 14648 23356 14724 23390
rect 14641 23340 14724 23356
rect 14539 23318 14724 23340
rect 14539 23306 14614 23318
rect 14539 23272 14607 23306
rect 14648 23284 14724 23318
rect 14641 23272 14724 23284
rect 14539 23246 14724 23272
rect 14539 23238 14614 23246
rect 14539 23204 14607 23238
rect 14648 23212 14724 23246
rect 14641 23204 14724 23212
rect 14539 23174 14724 23204
rect 14539 23170 14614 23174
rect 14539 23136 14607 23170
rect 14648 23140 14724 23174
rect 14641 23136 14724 23140
rect 14539 23102 14724 23136
rect 14539 23068 14607 23102
rect 14648 23068 14724 23102
rect 14539 23034 14724 23068
rect 14539 23000 14607 23034
rect 14641 23030 14724 23034
rect 14539 22996 14614 23000
rect 14648 22996 14724 23030
rect 14539 22966 14724 22996
rect 14539 22932 14607 22966
rect 14641 22958 14724 22966
rect 14539 22924 14614 22932
rect 14648 22924 14724 22958
rect 14539 22898 14724 22924
rect 14539 22864 14607 22898
rect 14641 22886 14724 22898
rect 14539 22852 14614 22864
rect 14648 22852 14724 22886
rect 14539 22830 14724 22852
rect 14539 22796 14607 22830
rect 14641 22814 14724 22830
rect 14539 22780 14614 22796
rect 14648 22780 14724 22814
rect 14539 22762 14724 22780
rect 14539 22728 14607 22762
rect 14641 22742 14724 22762
rect 14539 22708 14614 22728
rect 14648 22708 14724 22742
rect 14539 22694 14724 22708
rect 14539 22660 14607 22694
rect 14641 22670 14724 22694
rect 14539 22636 14614 22660
rect 14648 22636 14724 22670
rect 14539 22626 14724 22636
rect 14539 22592 14607 22626
rect 14641 22598 14724 22626
rect 14539 22564 14614 22592
rect 14648 22564 14724 22598
rect 14539 22558 14724 22564
rect 14539 22524 14607 22558
rect 14641 22526 14724 22558
rect 14539 22492 14614 22524
rect 14648 22492 14724 22526
rect 14539 22490 14724 22492
rect 14539 22456 14607 22490
rect 14641 22456 14724 22490
rect 14539 22454 14724 22456
rect 14539 22422 14614 22454
rect 14539 22388 14607 22422
rect 14648 22420 14724 22454
rect 14641 22388 14724 22420
rect 14539 22382 14724 22388
rect 14539 22354 14614 22382
rect 14539 22320 14607 22354
rect 14648 22348 14724 22382
rect 14641 22320 14724 22348
rect 14539 22310 14724 22320
rect 14539 22286 14614 22310
rect 14539 22252 14607 22286
rect 14648 22276 14724 22310
rect 14641 22252 14724 22276
rect 14539 22238 14724 22252
rect 14539 22218 14614 22238
rect 14539 22184 14607 22218
rect 14648 22204 14724 22238
rect 14641 22184 14724 22204
rect 14539 22166 14724 22184
rect 14539 22150 14614 22166
rect 14539 22116 14607 22150
rect 14648 22132 14724 22166
rect 14641 22116 14724 22132
rect 14539 22094 14724 22116
rect 14539 22082 14614 22094
rect 14539 22048 14607 22082
rect 14648 22060 14724 22094
rect 14641 22048 14724 22060
rect 14539 22022 14724 22048
rect 14539 22014 14614 22022
rect 14539 21980 14607 22014
rect 14648 21988 14724 22022
rect 14641 21980 14724 21988
rect 14539 21950 14724 21980
rect 14539 21946 14614 21950
rect 14539 21912 14607 21946
rect 14648 21916 14724 21950
rect 14641 21912 14724 21916
rect 14539 21878 14724 21912
rect 14539 21844 14607 21878
rect 14648 21844 14724 21878
rect 14539 21810 14724 21844
rect 14539 21776 14607 21810
rect 14641 21806 14724 21810
rect 14539 21772 14614 21776
rect 14648 21772 14724 21806
rect 14539 21742 14724 21772
rect 14539 21708 14607 21742
rect 14641 21734 14724 21742
rect 14539 21700 14614 21708
rect 14648 21700 14724 21734
rect 14539 21674 14724 21700
rect 14539 21640 14607 21674
rect 14641 21662 14724 21674
rect 14539 21628 14614 21640
rect 14648 21628 14724 21662
rect 14539 21606 14724 21628
rect 14539 21572 14607 21606
rect 14641 21590 14724 21606
rect 14539 21556 14614 21572
rect 14648 21556 14724 21590
rect 14539 21538 14724 21556
rect 14539 21504 14607 21538
rect 14641 21518 14724 21538
rect 14539 21484 14614 21504
rect 14648 21484 14724 21518
rect 14539 21470 14724 21484
rect 14539 21436 14607 21470
rect 14641 21446 14724 21470
rect 14539 21412 14614 21436
rect 14648 21412 14724 21446
rect 14539 21402 14724 21412
rect 14539 21368 14607 21402
rect 14641 21374 14724 21402
rect 14539 21340 14614 21368
rect 14648 21340 14724 21374
rect 14539 21334 14724 21340
rect 14539 21300 14607 21334
rect 14641 21302 14724 21334
rect 14539 21268 14614 21300
rect 14648 21268 14724 21302
rect 14539 21266 14724 21268
rect 14539 21232 14607 21266
rect 14641 21232 14724 21266
rect 14539 21230 14724 21232
rect 14539 21198 14614 21230
rect 14539 21164 14607 21198
rect 14648 21196 14724 21230
rect 14641 21164 14724 21196
rect 14539 21158 14724 21164
rect 14539 21130 14614 21158
rect 14539 21096 14607 21130
rect 14648 21124 14724 21158
rect 14641 21096 14724 21124
rect 14539 21086 14724 21096
rect 14539 21062 14614 21086
rect 14539 21028 14607 21062
rect 14648 21052 14724 21086
rect 14641 21028 14724 21052
rect 14539 21014 14724 21028
rect 14539 20994 14614 21014
rect 14539 20960 14607 20994
rect 14648 20980 14724 21014
rect 14641 20960 14724 20980
rect 14539 20942 14724 20960
rect 14539 20926 14614 20942
rect 14539 20892 14607 20926
rect 14648 20908 14724 20942
rect 14641 20892 14724 20908
rect 14539 20870 14724 20892
rect 14539 20858 14614 20870
rect 14539 20824 14607 20858
rect 14648 20836 14724 20870
rect 14641 20824 14724 20836
rect 14539 20798 14724 20824
rect 14539 20790 14614 20798
rect 14539 20756 14607 20790
rect 14648 20764 14724 20798
rect 14641 20756 14724 20764
rect 14539 20726 14724 20756
rect 14539 20722 14614 20726
rect 14539 20688 14607 20722
rect 14648 20692 14724 20726
rect 14641 20688 14724 20692
rect 14539 20654 14724 20688
rect 14539 20620 14607 20654
rect 14648 20620 14724 20654
rect 14539 20586 14724 20620
rect 14539 20552 14607 20586
rect 14641 20582 14724 20586
rect 14539 20548 14614 20552
rect 14648 20548 14724 20582
rect 14539 20518 14724 20548
rect 14539 20484 14607 20518
rect 14641 20510 14724 20518
rect 14539 20476 14614 20484
rect 14648 20476 14724 20510
rect 14539 20450 14724 20476
rect 14539 20416 14607 20450
rect 14641 20438 14724 20450
rect 14539 20404 14614 20416
rect 14648 20404 14724 20438
rect 14539 20382 14724 20404
rect 14539 20348 14607 20382
rect 14641 20366 14724 20382
rect 14539 20332 14614 20348
rect 14648 20332 14724 20366
rect 14539 20314 14724 20332
rect 14539 20280 14607 20314
rect 14641 20294 14724 20314
rect 14539 20260 14614 20280
rect 14648 20260 14724 20294
rect 14539 20246 14724 20260
rect 14539 20212 14607 20246
rect 14641 20222 14724 20246
rect 14539 20188 14614 20212
rect 14648 20188 14724 20222
rect 14539 20178 14724 20188
rect 14539 20144 14607 20178
rect 14641 20150 14724 20178
rect 14539 20116 14614 20144
rect 14648 20116 14724 20150
rect 14539 20110 14724 20116
rect 14539 20076 14607 20110
rect 14641 20078 14724 20110
rect 14539 20044 14614 20076
rect 14648 20044 14724 20078
rect 14539 20042 14724 20044
rect 14539 20008 14607 20042
rect 14641 20008 14724 20042
rect 14539 20006 14724 20008
rect 14539 19974 14614 20006
rect 14539 19940 14607 19974
rect 14648 19972 14724 20006
rect 14641 19940 14724 19972
rect 14539 19934 14724 19940
rect 14539 19906 14614 19934
rect 14539 19872 14607 19906
rect 14648 19900 14724 19934
rect 14641 19872 14724 19900
rect 14539 19862 14724 19872
rect 14539 19838 14614 19862
rect 14539 19804 14607 19838
rect 14648 19828 14724 19862
rect 14641 19804 14724 19828
rect 14539 19790 14724 19804
rect 14539 19770 14614 19790
rect 14539 19736 14607 19770
rect 14648 19756 14724 19790
rect 14641 19736 14724 19756
rect 14539 19718 14724 19736
rect 14539 19702 14614 19718
rect 14539 19668 14607 19702
rect 14648 19684 14724 19718
rect 14641 19668 14724 19684
rect 14539 19646 14724 19668
rect 14539 19634 14614 19646
rect 14539 19600 14607 19634
rect 14648 19612 14724 19646
rect 14641 19600 14724 19612
rect 14539 19574 14724 19600
rect 14539 19566 14614 19574
rect 14539 19532 14607 19566
rect 14648 19540 14724 19574
rect 14641 19532 14724 19540
rect 14539 19502 14724 19532
rect 14539 19498 14614 19502
rect 14539 19464 14607 19498
rect 14648 19468 14724 19502
rect 14641 19464 14724 19468
rect 14539 19430 14724 19464
rect 14539 19396 14607 19430
rect 14648 19396 14724 19430
rect 14539 19362 14724 19396
rect 14539 19328 14607 19362
rect 14641 19358 14724 19362
rect 14539 19324 14614 19328
rect 14648 19324 14724 19358
rect 14539 19294 14724 19324
rect 14539 19260 14607 19294
rect 14641 19286 14724 19294
rect 14539 19252 14614 19260
rect 14648 19252 14724 19286
rect 14539 19226 14724 19252
rect 14539 19192 14607 19226
rect 14641 19214 14724 19226
rect 14539 19180 14614 19192
rect 14648 19180 14724 19214
rect 14539 19158 14724 19180
rect 14539 19124 14607 19158
rect 14641 19142 14724 19158
rect 14539 19108 14614 19124
rect 14648 19108 14724 19142
rect 14539 19090 14724 19108
rect 14539 19056 14607 19090
rect 14641 19070 14724 19090
rect 14539 19036 14614 19056
rect 14648 19036 14724 19070
rect 14539 19022 14724 19036
rect 14539 18988 14607 19022
rect 14641 18998 14724 19022
rect 14539 18964 14614 18988
rect 14648 18964 14724 18998
rect 14539 18954 14724 18964
rect 14539 18920 14607 18954
rect 14641 18926 14724 18954
rect 14539 18892 14614 18920
rect 14648 18892 14724 18926
rect 14539 18886 14724 18892
rect 14539 18852 14607 18886
rect 14641 18854 14724 18886
rect 14539 18820 14614 18852
rect 14648 18820 14724 18854
rect 14539 18818 14724 18820
rect 14539 18784 14607 18818
rect 14641 18784 14724 18818
rect 14539 18782 14724 18784
rect 14539 18750 14614 18782
rect 14539 18716 14607 18750
rect 14648 18748 14724 18782
rect 14641 18716 14724 18748
rect 14539 18710 14724 18716
rect 14539 18682 14614 18710
rect 14539 18648 14607 18682
rect 14648 18676 14724 18710
rect 14641 18648 14724 18676
rect 14539 18638 14724 18648
rect 14539 18614 14614 18638
rect 14539 18580 14607 18614
rect 14648 18604 14724 18638
rect 14641 18580 14724 18604
rect 14539 18566 14724 18580
rect 14539 18546 14614 18566
rect 14539 18512 14607 18546
rect 14648 18532 14724 18566
rect 14641 18512 14724 18532
rect 14539 18494 14724 18512
rect 14539 18478 14614 18494
rect 14539 18444 14607 18478
rect 14648 18460 14724 18494
rect 14641 18444 14724 18460
rect 14539 18422 14724 18444
rect 14539 18410 14614 18422
rect 14539 18376 14607 18410
rect 14648 18388 14724 18422
rect 14641 18376 14724 18388
rect 14539 18350 14724 18376
rect 14539 18342 14614 18350
rect 14539 18308 14607 18342
rect 14648 18316 14724 18350
rect 14641 18308 14724 18316
rect 14539 18278 14724 18308
rect 14539 18274 14614 18278
rect 14539 18240 14607 18274
rect 14648 18244 14724 18278
rect 14641 18240 14724 18244
rect 14539 18206 14724 18240
rect 14539 18172 14607 18206
rect 14648 18172 14724 18206
rect 14539 18138 14724 18172
rect 14539 18104 14607 18138
rect 14641 18134 14724 18138
rect 14539 18100 14614 18104
rect 14648 18100 14724 18134
rect 14539 18070 14724 18100
rect 14539 18036 14607 18070
rect 14641 18062 14724 18070
rect 14539 18028 14614 18036
rect 14648 18028 14724 18062
rect 14539 18002 14724 18028
rect 14539 17968 14607 18002
rect 14641 17990 14724 18002
rect 14539 17956 14614 17968
rect 14648 17956 14724 17990
rect 14539 17934 14724 17956
rect 14539 17900 14607 17934
rect 14641 17918 14724 17934
rect 14539 17884 14614 17900
rect 14648 17884 14724 17918
rect 14539 17866 14724 17884
rect 14539 17832 14607 17866
rect 14641 17846 14724 17866
rect 14539 17812 14614 17832
rect 14648 17812 14724 17846
rect 14539 17798 14724 17812
rect 14539 17764 14607 17798
rect 14641 17774 14724 17798
rect 14539 17740 14614 17764
rect 14648 17740 14724 17774
rect 14539 17730 14724 17740
rect 14539 17696 14607 17730
rect 14641 17702 14724 17730
rect 14539 17668 14614 17696
rect 14648 17668 14724 17702
rect 14539 17662 14724 17668
rect 14539 17628 14607 17662
rect 14641 17630 14724 17662
rect 14539 17596 14614 17628
rect 14648 17596 14724 17630
rect 14539 17594 14724 17596
rect 14539 17560 14607 17594
rect 14641 17560 14724 17594
rect 14539 17558 14724 17560
rect 14539 17526 14614 17558
rect 14539 17492 14607 17526
rect 14648 17524 14724 17558
rect 14641 17492 14724 17524
rect 14539 17486 14724 17492
rect 14539 17458 14614 17486
rect 14539 17424 14607 17458
rect 14648 17452 14724 17486
rect 14641 17424 14724 17452
rect 14539 17414 14724 17424
rect 14539 17390 14614 17414
rect 14539 17356 14607 17390
rect 14648 17380 14724 17414
rect 14641 17356 14724 17380
rect 14539 17342 14724 17356
rect 14539 17322 14614 17342
rect 14539 17288 14607 17322
rect 14648 17308 14724 17342
rect 14641 17288 14724 17308
rect 14539 17270 14724 17288
rect 14539 17254 14614 17270
rect 14539 17220 14607 17254
rect 14648 17236 14724 17270
rect 14641 17220 14724 17236
rect 14539 17198 14724 17220
rect 14539 17186 14614 17198
rect 14539 17152 14607 17186
rect 14648 17164 14724 17198
rect 14641 17152 14724 17164
rect 14539 17126 14724 17152
rect 14539 17118 14614 17126
rect 14539 17084 14607 17118
rect 14648 17092 14724 17126
rect 14641 17084 14724 17092
rect 14539 17054 14724 17084
rect 14539 17050 14614 17054
rect 14539 17016 14607 17050
rect 14648 17020 14724 17054
rect 14641 17016 14724 17020
rect 14539 16982 14724 17016
rect 14539 16948 14607 16982
rect 14648 16948 14724 16982
rect 14539 16914 14724 16948
rect 14539 16880 14607 16914
rect 14641 16910 14724 16914
rect 14539 16876 14614 16880
rect 14648 16876 14724 16910
rect 14539 16846 14724 16876
rect 14539 16812 14607 16846
rect 14641 16838 14724 16846
rect 14539 16804 14614 16812
rect 14648 16804 14724 16838
rect 14539 16778 14724 16804
rect 14539 16744 14607 16778
rect 14641 16766 14724 16778
rect 14539 16732 14614 16744
rect 14648 16732 14724 16766
rect 14539 16710 14724 16732
rect 14539 16676 14607 16710
rect 14641 16694 14724 16710
rect 14539 16660 14614 16676
rect 14648 16660 14724 16694
rect 14539 16642 14724 16660
rect 14539 16608 14607 16642
rect 14641 16622 14724 16642
rect 14539 16588 14614 16608
rect 14648 16588 14724 16622
rect 14539 16574 14724 16588
rect 14539 16540 14607 16574
rect 14641 16550 14724 16574
rect 14539 16516 14614 16540
rect 14648 16516 14724 16550
rect 14539 16506 14724 16516
rect 14539 16472 14607 16506
rect 14641 16478 14724 16506
rect 14539 16444 14614 16472
rect 14648 16444 14724 16478
rect 14539 16438 14724 16444
rect 14539 16404 14607 16438
rect 14641 16406 14724 16438
rect 14539 16372 14614 16404
rect 14648 16372 14724 16406
rect 14539 16370 14724 16372
rect 14539 16336 14607 16370
rect 14641 16336 14724 16370
rect 14539 16334 14724 16336
rect 14539 16302 14614 16334
rect 14539 16268 14607 16302
rect 14648 16300 14724 16334
rect 14641 16268 14724 16300
rect 14539 16262 14724 16268
rect 14539 16234 14614 16262
rect 14539 16200 14607 16234
rect 14648 16228 14724 16262
rect 14641 16200 14724 16228
rect 14539 16190 14724 16200
rect 14539 16166 14614 16190
rect 14539 16132 14607 16166
rect 14648 16156 14724 16190
rect 14641 16132 14724 16156
rect 14539 16118 14724 16132
rect 14539 16098 14614 16118
rect 14539 16064 14607 16098
rect 14648 16084 14724 16118
rect 14641 16064 14724 16084
rect 14539 16046 14724 16064
rect 14539 16030 14614 16046
rect 14539 15996 14607 16030
rect 14648 16012 14724 16046
rect 14641 15996 14724 16012
rect 14539 15974 14724 15996
rect 14539 15962 14614 15974
rect 14539 15928 14607 15962
rect 14648 15940 14724 15974
rect 14641 15928 14724 15940
rect 14539 15902 14724 15928
rect 14539 15894 14614 15902
rect 14539 15860 14607 15894
rect 14648 15868 14724 15902
rect 14641 15860 14724 15868
rect 14539 15830 14724 15860
rect 14539 15826 14614 15830
rect 14539 15792 14607 15826
rect 14648 15796 14724 15830
rect 14641 15792 14724 15796
rect 14539 15758 14724 15792
rect 14539 15724 14607 15758
rect 14648 15724 14724 15758
rect 14539 15690 14724 15724
rect 14539 15656 14607 15690
rect 14641 15686 14724 15690
rect 14539 15652 14614 15656
rect 14648 15652 14724 15686
rect 14539 15622 14724 15652
rect 14539 15588 14607 15622
rect 14641 15614 14724 15622
rect 14539 15580 14614 15588
rect 14648 15580 14724 15614
rect 14539 15554 14724 15580
rect 14539 15520 14607 15554
rect 14641 15542 14724 15554
rect 14539 15508 14614 15520
rect 14648 15508 14724 15542
rect 14539 15486 14724 15508
rect 14539 15452 14607 15486
rect 14641 15470 14724 15486
rect 14539 15436 14614 15452
rect 14648 15436 14724 15470
rect 14539 15418 14724 15436
rect 14539 15384 14607 15418
rect 14641 15398 14724 15418
rect 14539 15364 14614 15384
rect 14648 15364 14724 15398
rect 14539 15350 14724 15364
rect 14539 15316 14607 15350
rect 14641 15326 14724 15350
rect 14539 15292 14614 15316
rect 14648 15292 14724 15326
rect 14539 15282 14724 15292
rect 14539 15248 14607 15282
rect 14641 15254 14724 15282
rect 14539 15220 14614 15248
rect 14648 15220 14724 15254
rect 14539 15214 14724 15220
rect 14539 15180 14607 15214
rect 14641 15182 14724 15214
rect 14539 15148 14614 15180
rect 14648 15148 14724 15182
rect 14539 15146 14724 15148
rect 14539 15112 14607 15146
rect 14641 15112 14724 15146
rect 14539 15110 14724 15112
rect 14539 15078 14614 15110
rect 14539 15044 14607 15078
rect 14648 15076 14724 15110
rect 14641 15044 14724 15076
rect 14539 15038 14724 15044
rect 14539 15010 14614 15038
rect 14539 14976 14607 15010
rect 14648 15004 14724 15038
rect 14641 14976 14724 15004
rect 14539 14966 14724 14976
rect 14539 14942 14614 14966
rect 14539 14908 14607 14942
rect 14648 14932 14724 14966
rect 14641 14908 14724 14932
rect 14539 14894 14724 14908
rect 14539 14874 14614 14894
rect 14539 14840 14607 14874
rect 14648 14860 14724 14894
rect 14641 14840 14724 14860
rect 14539 14822 14724 14840
rect 14539 14806 14614 14822
rect 14539 14772 14607 14806
rect 14648 14788 14724 14822
rect 14641 14772 14724 14788
rect 14539 14750 14724 14772
rect 14539 14738 14614 14750
rect 882 14710 2070 14711
rect 12882 14710 14070 14711
rect 245 14681 430 14698
rect 245 14664 320 14681
rect 245 14630 312 14664
rect 354 14647 430 14681
rect 346 14630 430 14647
rect 245 14596 430 14630
rect 245 14562 312 14596
rect 346 14562 430 14596
rect 245 14528 430 14562
rect 14539 14704 14607 14738
rect 14648 14716 14724 14750
rect 14641 14704 14724 14716
rect 14539 14678 14724 14704
rect 14539 14670 14614 14678
rect 14539 14636 14607 14670
rect 14648 14644 14724 14678
rect 14641 14636 14724 14644
rect 14539 14602 14724 14636
rect 14539 14568 14607 14602
rect 14641 14568 14724 14602
rect 14539 14528 14724 14568
rect 245 14452 14724 14528
rect 245 14418 320 14452
rect 354 14451 610 14452
rect 644 14451 2311 14452
rect 2345 14451 2383 14452
rect 2417 14451 2455 14452
rect 2489 14451 2527 14452
rect 2561 14451 2599 14452
rect 2633 14451 2671 14452
rect 2705 14451 2743 14452
rect 2777 14451 2815 14452
rect 2849 14451 2887 14452
rect 2921 14451 2959 14452
rect 2993 14451 3031 14452
rect 3065 14451 3103 14452
rect 3137 14451 3175 14452
rect 3209 14451 3247 14452
rect 3281 14451 3319 14452
rect 3353 14451 3391 14452
rect 3425 14451 3463 14452
rect 3497 14451 3535 14452
rect 3569 14451 3607 14452
rect 3641 14451 3679 14452
rect 3713 14451 3751 14452
rect 3785 14451 3823 14452
rect 3857 14451 3895 14452
rect 3929 14451 3967 14452
rect 4001 14451 4039 14452
rect 4073 14451 4111 14452
rect 4145 14451 4183 14452
rect 4217 14451 4255 14452
rect 4289 14451 4327 14452
rect 4361 14451 4399 14452
rect 4433 14451 4471 14452
rect 4505 14451 4543 14452
rect 4577 14451 4615 14452
rect 4649 14451 4687 14452
rect 4721 14451 4759 14452
rect 4793 14451 4831 14452
rect 4865 14451 4903 14452
rect 4937 14451 4975 14452
rect 5009 14451 5047 14452
rect 5081 14451 5119 14452
rect 5153 14451 5191 14452
rect 5225 14451 5263 14452
rect 5297 14451 5335 14452
rect 5369 14451 5407 14452
rect 5441 14451 5479 14452
rect 5513 14451 5551 14452
rect 5585 14451 5623 14452
rect 5657 14451 5695 14452
rect 5729 14451 5767 14452
rect 5801 14451 5839 14452
rect 5873 14451 5911 14452
rect 5945 14451 5983 14452
rect 6017 14451 6055 14452
rect 6089 14451 6127 14452
rect 6161 14451 6199 14452
rect 6233 14451 6271 14452
rect 6305 14451 6343 14452
rect 6377 14451 6415 14452
rect 6449 14451 6487 14452
rect 6521 14451 6559 14452
rect 6593 14451 6631 14452
rect 6665 14451 6703 14452
rect 6737 14451 6775 14452
rect 6809 14451 6847 14452
rect 6881 14451 6919 14452
rect 6953 14451 6991 14452
rect 7025 14451 7063 14452
rect 7097 14451 7135 14452
rect 7169 14451 7207 14452
rect 7241 14451 7279 14452
rect 7313 14451 7351 14452
rect 7385 14451 7423 14452
rect 7457 14451 7495 14452
rect 7529 14451 7567 14452
rect 7601 14451 7639 14452
rect 7673 14451 7711 14452
rect 7745 14451 7783 14452
rect 7817 14451 7855 14452
rect 7889 14451 7927 14452
rect 7961 14451 7999 14452
rect 8033 14451 8071 14452
rect 8105 14451 8143 14452
rect 8177 14451 8215 14452
rect 8249 14451 8287 14452
rect 8321 14451 8359 14452
rect 8393 14451 8431 14452
rect 8465 14451 8503 14452
rect 8537 14451 8575 14452
rect 8609 14451 8647 14452
rect 8681 14451 8719 14452
rect 8753 14451 8791 14452
rect 8825 14451 8863 14452
rect 8897 14451 8935 14452
rect 8969 14451 9007 14452
rect 9041 14451 9079 14452
rect 9113 14451 9151 14452
rect 9185 14451 9223 14452
rect 9257 14451 9295 14452
rect 9329 14451 9367 14452
rect 9401 14451 9439 14452
rect 9473 14451 9511 14452
rect 9545 14451 9583 14452
rect 9617 14451 9655 14452
rect 9689 14451 9727 14452
rect 9761 14451 9799 14452
rect 9833 14451 9871 14452
rect 9905 14451 9943 14452
rect 9977 14451 10015 14452
rect 10049 14451 10087 14452
rect 10121 14451 10159 14452
rect 10193 14451 10231 14452
rect 10265 14451 10303 14452
rect 10337 14451 10375 14452
rect 10409 14451 10447 14452
rect 10481 14451 10519 14452
rect 10553 14451 10591 14452
rect 10625 14451 10663 14452
rect 10697 14451 10735 14452
rect 10769 14451 10807 14452
rect 10841 14451 10879 14452
rect 10913 14451 10951 14452
rect 10985 14451 11023 14452
rect 11057 14451 11095 14452
rect 11129 14451 11167 14452
rect 11201 14451 11239 14452
rect 11273 14451 11311 14452
rect 11345 14451 11383 14452
rect 11417 14451 11455 14452
rect 11489 14451 11527 14452
rect 11561 14451 11599 14452
rect 11633 14451 11671 14452
rect 11705 14451 11743 14452
rect 11777 14451 11815 14452
rect 11849 14451 11887 14452
rect 11921 14451 11959 14452
rect 11993 14451 12031 14452
rect 12065 14451 12103 14452
rect 12137 14451 12175 14452
rect 12209 14451 12247 14452
rect 12281 14451 12319 14452
rect 12353 14451 12391 14452
rect 12425 14451 12463 14452
rect 12497 14451 12535 14452
rect 12569 14451 12607 14452
rect 12641 14451 14314 14452
rect 354 14418 476 14451
rect 245 14417 476 14418
rect 510 14417 544 14451
rect 578 14418 610 14451
rect 578 14417 612 14418
rect 646 14417 680 14451
rect 714 14417 748 14451
rect 782 14417 816 14451
rect 850 14417 884 14451
rect 918 14417 952 14451
rect 986 14417 1020 14451
rect 1054 14417 1088 14451
rect 1122 14417 1156 14451
rect 1190 14417 1224 14451
rect 1258 14417 1292 14451
rect 1326 14417 1360 14451
rect 1394 14417 1428 14451
rect 1462 14417 1496 14451
rect 1530 14417 1564 14451
rect 1598 14417 1632 14451
rect 1666 14417 1700 14451
rect 1734 14417 1768 14451
rect 1802 14417 1836 14451
rect 1870 14417 1904 14451
rect 1938 14417 1972 14451
rect 2006 14417 2040 14451
rect 2074 14417 2108 14451
rect 2142 14417 2176 14451
rect 2210 14417 2244 14451
rect 2278 14418 2311 14451
rect 2278 14417 2312 14418
rect 2346 14417 2380 14451
rect 2417 14418 2448 14451
rect 2489 14418 2516 14451
rect 2561 14418 2584 14451
rect 2633 14418 2652 14451
rect 2705 14418 2720 14451
rect 2777 14418 2788 14451
rect 2849 14418 2856 14451
rect 2921 14418 2924 14451
rect 2414 14417 2448 14418
rect 2482 14417 2516 14418
rect 2550 14417 2584 14418
rect 2618 14417 2652 14418
rect 2686 14417 2720 14418
rect 2754 14417 2788 14418
rect 2822 14417 2856 14418
rect 2890 14417 2924 14418
rect 2958 14418 2959 14451
rect 3026 14418 3031 14451
rect 3094 14418 3103 14451
rect 3162 14418 3175 14451
rect 3230 14418 3247 14451
rect 3298 14418 3319 14451
rect 3366 14418 3391 14451
rect 3434 14418 3463 14451
rect 3502 14418 3535 14451
rect 2958 14417 2992 14418
rect 3026 14417 3060 14418
rect 3094 14417 3128 14418
rect 3162 14417 3196 14418
rect 3230 14417 3264 14418
rect 3298 14417 3332 14418
rect 3366 14417 3400 14418
rect 3434 14417 3468 14418
rect 3502 14417 3536 14418
rect 3570 14417 3604 14451
rect 3641 14418 3672 14451
rect 3713 14418 3740 14451
rect 3785 14418 3808 14451
rect 3857 14418 3876 14451
rect 3929 14418 3944 14451
rect 4001 14418 4012 14451
rect 4073 14418 4080 14451
rect 4145 14418 4148 14451
rect 3638 14417 3672 14418
rect 3706 14417 3740 14418
rect 3774 14417 3808 14418
rect 3842 14417 3876 14418
rect 3910 14417 3944 14418
rect 3978 14417 4012 14418
rect 4046 14417 4080 14418
rect 4114 14417 4148 14418
rect 4182 14418 4183 14451
rect 4250 14418 4255 14451
rect 4318 14418 4327 14451
rect 4386 14418 4399 14451
rect 4454 14418 4471 14451
rect 4522 14418 4543 14451
rect 4590 14418 4615 14451
rect 4658 14418 4687 14451
rect 4726 14418 4759 14451
rect 4182 14417 4216 14418
rect 4250 14417 4284 14418
rect 4318 14417 4352 14418
rect 4386 14417 4420 14418
rect 4454 14417 4488 14418
rect 4522 14417 4556 14418
rect 4590 14417 4624 14418
rect 4658 14417 4692 14418
rect 4726 14417 4760 14418
rect 4794 14417 4828 14451
rect 4865 14418 4896 14451
rect 4937 14418 4964 14451
rect 5009 14418 5032 14451
rect 5081 14418 5100 14451
rect 5153 14418 5168 14451
rect 5225 14418 5236 14451
rect 5297 14418 5304 14451
rect 5369 14418 5372 14451
rect 4862 14417 4896 14418
rect 4930 14417 4964 14418
rect 4998 14417 5032 14418
rect 5066 14417 5100 14418
rect 5134 14417 5168 14418
rect 5202 14417 5236 14418
rect 5270 14417 5304 14418
rect 5338 14417 5372 14418
rect 5406 14418 5407 14451
rect 5474 14418 5479 14451
rect 5542 14418 5551 14451
rect 5610 14418 5623 14451
rect 5678 14418 5695 14451
rect 5746 14418 5767 14451
rect 5814 14418 5839 14451
rect 5882 14418 5911 14451
rect 5950 14418 5983 14451
rect 5406 14417 5440 14418
rect 5474 14417 5508 14418
rect 5542 14417 5576 14418
rect 5610 14417 5644 14418
rect 5678 14417 5712 14418
rect 5746 14417 5780 14418
rect 5814 14417 5848 14418
rect 5882 14417 5916 14418
rect 5950 14417 5984 14418
rect 6018 14417 6052 14451
rect 6089 14418 6120 14451
rect 6161 14418 6188 14451
rect 6233 14418 6256 14451
rect 6305 14418 6324 14451
rect 6377 14418 6392 14451
rect 6449 14418 6460 14451
rect 6521 14418 6528 14451
rect 6593 14418 6596 14451
rect 6086 14417 6120 14418
rect 6154 14417 6188 14418
rect 6222 14417 6256 14418
rect 6290 14417 6324 14418
rect 6358 14417 6392 14418
rect 6426 14417 6460 14418
rect 6494 14417 6528 14418
rect 6562 14417 6596 14418
rect 6630 14418 6631 14451
rect 6698 14418 6703 14451
rect 6766 14418 6775 14451
rect 6834 14418 6847 14451
rect 6902 14418 6919 14451
rect 6970 14418 6991 14451
rect 7038 14418 7063 14451
rect 7106 14418 7135 14451
rect 7174 14418 7207 14451
rect 6630 14417 6664 14418
rect 6698 14417 6732 14418
rect 6766 14417 6800 14418
rect 6834 14417 6868 14418
rect 6902 14417 6936 14418
rect 6970 14417 7004 14418
rect 7038 14417 7072 14418
rect 7106 14417 7140 14418
rect 7174 14417 7208 14418
rect 7242 14417 7276 14451
rect 7313 14418 7344 14451
rect 7385 14418 7412 14451
rect 7457 14418 7480 14451
rect 7529 14418 7548 14451
rect 7601 14418 7616 14451
rect 7673 14418 7684 14451
rect 7745 14418 7752 14451
rect 7817 14418 7820 14451
rect 7310 14417 7344 14418
rect 7378 14417 7412 14418
rect 7446 14417 7480 14418
rect 7514 14417 7548 14418
rect 7582 14417 7616 14418
rect 7650 14417 7684 14418
rect 7718 14417 7752 14418
rect 7786 14417 7820 14418
rect 7854 14418 7855 14451
rect 7922 14418 7927 14451
rect 7990 14418 7999 14451
rect 8058 14418 8071 14451
rect 8126 14418 8143 14451
rect 8194 14418 8215 14451
rect 8262 14418 8287 14451
rect 8330 14418 8359 14451
rect 8398 14418 8431 14451
rect 7854 14417 7888 14418
rect 7922 14417 7956 14418
rect 7990 14417 8024 14418
rect 8058 14417 8092 14418
rect 8126 14417 8160 14418
rect 8194 14417 8228 14418
rect 8262 14417 8296 14418
rect 8330 14417 8364 14418
rect 8398 14417 8432 14418
rect 8466 14417 8500 14451
rect 8537 14418 8568 14451
rect 8609 14418 8636 14451
rect 8681 14418 8704 14451
rect 8753 14418 8772 14451
rect 8825 14418 8840 14451
rect 8897 14418 8908 14451
rect 8969 14418 8976 14451
rect 9041 14418 9044 14451
rect 8534 14417 8568 14418
rect 8602 14417 8636 14418
rect 8670 14417 8704 14418
rect 8738 14417 8772 14418
rect 8806 14417 8840 14418
rect 8874 14417 8908 14418
rect 8942 14417 8976 14418
rect 9010 14417 9044 14418
rect 9078 14418 9079 14451
rect 9146 14418 9151 14451
rect 9214 14418 9223 14451
rect 9282 14418 9295 14451
rect 9350 14418 9367 14451
rect 9418 14418 9439 14451
rect 9486 14418 9511 14451
rect 9554 14418 9583 14451
rect 9622 14418 9655 14451
rect 9078 14417 9112 14418
rect 9146 14417 9180 14418
rect 9214 14417 9248 14418
rect 9282 14417 9316 14418
rect 9350 14417 9384 14418
rect 9418 14417 9452 14418
rect 9486 14417 9520 14418
rect 9554 14417 9588 14418
rect 9622 14417 9656 14418
rect 9690 14417 9724 14451
rect 9761 14418 9792 14451
rect 9833 14418 9860 14451
rect 9905 14418 9928 14451
rect 9977 14418 9996 14451
rect 10049 14418 10064 14451
rect 10121 14418 10132 14451
rect 10193 14418 10200 14451
rect 10265 14418 10268 14451
rect 9758 14417 9792 14418
rect 9826 14417 9860 14418
rect 9894 14417 9928 14418
rect 9962 14417 9996 14418
rect 10030 14417 10064 14418
rect 10098 14417 10132 14418
rect 10166 14417 10200 14418
rect 10234 14417 10268 14418
rect 10302 14418 10303 14451
rect 10370 14418 10375 14451
rect 10438 14418 10447 14451
rect 10506 14418 10519 14451
rect 10574 14418 10591 14451
rect 10642 14418 10663 14451
rect 10710 14418 10735 14451
rect 10778 14418 10807 14451
rect 10846 14418 10879 14451
rect 10302 14417 10336 14418
rect 10370 14417 10404 14418
rect 10438 14417 10472 14418
rect 10506 14417 10540 14418
rect 10574 14417 10608 14418
rect 10642 14417 10676 14418
rect 10710 14417 10744 14418
rect 10778 14417 10812 14418
rect 10846 14417 10880 14418
rect 10914 14417 10948 14451
rect 10985 14418 11016 14451
rect 11057 14418 11084 14451
rect 11129 14418 11152 14451
rect 11201 14418 11220 14451
rect 11273 14418 11288 14451
rect 11345 14418 11356 14451
rect 11417 14418 11424 14451
rect 11489 14418 11492 14451
rect 10982 14417 11016 14418
rect 11050 14417 11084 14418
rect 11118 14417 11152 14418
rect 11186 14417 11220 14418
rect 11254 14417 11288 14418
rect 11322 14417 11356 14418
rect 11390 14417 11424 14418
rect 11458 14417 11492 14418
rect 11526 14418 11527 14451
rect 11594 14418 11599 14451
rect 11662 14418 11671 14451
rect 11730 14418 11743 14451
rect 11798 14418 11815 14451
rect 11866 14418 11887 14451
rect 11934 14418 11959 14451
rect 12002 14418 12031 14451
rect 12070 14418 12103 14451
rect 11526 14417 11560 14418
rect 11594 14417 11628 14418
rect 11662 14417 11696 14418
rect 11730 14417 11764 14418
rect 11798 14417 11832 14418
rect 11866 14417 11900 14418
rect 11934 14417 11968 14418
rect 12002 14417 12036 14418
rect 12070 14417 12104 14418
rect 12138 14417 12172 14451
rect 12209 14418 12240 14451
rect 12281 14418 12308 14451
rect 12353 14418 12376 14451
rect 12425 14418 12444 14451
rect 12497 14418 12512 14451
rect 12569 14418 12580 14451
rect 12641 14418 12648 14451
rect 12206 14417 12240 14418
rect 12274 14417 12308 14418
rect 12342 14417 12376 14418
rect 12410 14417 12444 14418
rect 12478 14417 12512 14418
rect 12546 14417 12580 14418
rect 12614 14417 12648 14418
rect 12682 14417 12716 14451
rect 12750 14417 12784 14451
rect 12818 14417 12852 14451
rect 12886 14417 12920 14451
rect 12954 14417 12988 14451
rect 13022 14417 13056 14451
rect 13090 14417 13124 14451
rect 13158 14417 13192 14451
rect 13226 14417 13260 14451
rect 13294 14417 13328 14451
rect 13362 14417 13396 14451
rect 13430 14417 13464 14451
rect 13498 14417 13532 14451
rect 13566 14417 13600 14451
rect 13634 14417 13668 14451
rect 13702 14417 13736 14451
rect 13770 14417 13804 14451
rect 13838 14417 13872 14451
rect 13906 14417 13940 14451
rect 13974 14417 14008 14451
rect 14042 14417 14076 14451
rect 14110 14417 14144 14451
rect 14178 14417 14212 14451
rect 14246 14417 14280 14451
rect 14348 14451 14614 14452
rect 14314 14417 14348 14418
rect 14382 14417 14416 14451
rect 14450 14417 14484 14451
rect 14518 14418 14614 14451
rect 14648 14418 14724 14452
rect 14518 14417 14724 14418
rect 245 14343 14724 14417
<< viali >>
rect 320 36500 354 36534
rect 14614 36499 14648 36533
rect 556 36497 590 36498
rect 628 36497 662 36498
rect 700 36497 734 36498
rect 772 36497 806 36498
rect 844 36497 878 36498
rect 916 36497 950 36498
rect 988 36497 1022 36498
rect 1060 36497 1094 36498
rect 1132 36497 1166 36498
rect 1204 36497 1238 36498
rect 1276 36497 1310 36498
rect 1348 36497 1382 36498
rect 1420 36497 1454 36498
rect 1492 36497 1526 36498
rect 1564 36497 1598 36498
rect 1636 36497 1670 36498
rect 1708 36497 1742 36498
rect 1780 36497 1814 36498
rect 1852 36497 1886 36498
rect 1924 36497 1958 36498
rect 1996 36497 2030 36498
rect 2068 36497 2102 36498
rect 2140 36497 2174 36498
rect 2212 36497 2246 36498
rect 2284 36497 2318 36498
rect 2356 36497 2390 36498
rect 2428 36497 2462 36498
rect 2500 36497 2534 36498
rect 2572 36497 2606 36498
rect 2644 36497 2678 36498
rect 2716 36497 2750 36498
rect 2788 36497 2822 36498
rect 2860 36497 2894 36498
rect 2932 36497 2966 36498
rect 3004 36497 3038 36498
rect 3076 36497 3110 36498
rect 3148 36497 3182 36498
rect 3220 36497 3254 36498
rect 3292 36497 3326 36498
rect 3364 36497 3398 36498
rect 3436 36497 3470 36498
rect 3508 36497 3542 36498
rect 3580 36497 3614 36498
rect 3652 36497 3686 36498
rect 3724 36497 3758 36498
rect 3796 36497 3830 36498
rect 3868 36497 3902 36498
rect 3940 36497 3974 36498
rect 4012 36497 4046 36498
rect 4084 36497 4118 36498
rect 4156 36497 4190 36498
rect 4228 36497 4262 36498
rect 4300 36497 4334 36498
rect 4372 36497 4406 36498
rect 4444 36497 4478 36498
rect 4516 36497 4550 36498
rect 4588 36497 4622 36498
rect 4660 36497 4694 36498
rect 4732 36497 4766 36498
rect 4804 36497 4838 36498
rect 4876 36497 4910 36498
rect 4948 36497 4982 36498
rect 5020 36497 5054 36498
rect 5092 36497 5126 36498
rect 5164 36497 5198 36498
rect 5236 36497 5270 36498
rect 5308 36497 5342 36498
rect 5380 36497 5414 36498
rect 5452 36497 5486 36498
rect 5524 36497 5558 36498
rect 5596 36497 5630 36498
rect 5668 36497 5702 36498
rect 5740 36497 5774 36498
rect 5812 36497 5846 36498
rect 5884 36497 5918 36498
rect 5956 36497 5990 36498
rect 6028 36497 6062 36498
rect 6100 36497 6134 36498
rect 6172 36497 6206 36498
rect 6244 36497 6278 36498
rect 6316 36497 6350 36498
rect 6388 36497 6422 36498
rect 6460 36497 6494 36498
rect 6532 36497 6566 36498
rect 6604 36497 6638 36498
rect 6676 36497 6710 36498
rect 6748 36497 6782 36498
rect 6820 36497 6854 36498
rect 6892 36497 6926 36498
rect 6964 36497 6998 36498
rect 7036 36497 7070 36498
rect 7108 36497 7142 36498
rect 7180 36497 7214 36498
rect 7252 36497 7286 36498
rect 7324 36497 7358 36498
rect 7396 36497 7430 36498
rect 7468 36497 7502 36498
rect 7540 36497 7574 36498
rect 7612 36497 7646 36498
rect 7684 36497 7718 36498
rect 7756 36497 7790 36498
rect 7828 36497 7862 36498
rect 7900 36497 7934 36498
rect 7972 36497 8006 36498
rect 8044 36497 8078 36498
rect 8116 36497 8150 36498
rect 8188 36497 8222 36498
rect 8260 36497 8294 36498
rect 8332 36497 8366 36498
rect 8404 36497 8438 36498
rect 8476 36497 8510 36498
rect 8548 36497 8582 36498
rect 8620 36497 8654 36498
rect 8692 36497 8726 36498
rect 8764 36497 8798 36498
rect 8836 36497 8870 36498
rect 8908 36497 8942 36498
rect 8980 36497 9014 36498
rect 9052 36497 9086 36498
rect 9124 36497 9158 36498
rect 9196 36497 9230 36498
rect 9268 36497 9302 36498
rect 9340 36497 9374 36498
rect 9412 36497 9446 36498
rect 9484 36497 9518 36498
rect 9556 36497 9590 36498
rect 9628 36497 9662 36498
rect 9700 36497 9734 36498
rect 9772 36497 9806 36498
rect 9844 36497 9878 36498
rect 9916 36497 9950 36498
rect 9988 36497 10022 36498
rect 10060 36497 10094 36498
rect 10132 36497 10166 36498
rect 10204 36497 10238 36498
rect 10276 36497 10310 36498
rect 10348 36497 10382 36498
rect 10420 36497 10454 36498
rect 10492 36497 10526 36498
rect 10564 36497 10598 36498
rect 10636 36497 10670 36498
rect 10708 36497 10742 36498
rect 10780 36497 10814 36498
rect 10852 36497 10886 36498
rect 10924 36497 10958 36498
rect 10996 36497 11030 36498
rect 11068 36497 11102 36498
rect 11140 36497 11174 36498
rect 11212 36497 11246 36498
rect 11284 36497 11318 36498
rect 11356 36497 11390 36498
rect 11428 36497 11462 36498
rect 11500 36497 11534 36498
rect 11572 36497 11606 36498
rect 11644 36497 11678 36498
rect 11716 36497 11750 36498
rect 11788 36497 11822 36498
rect 11860 36497 11894 36498
rect 11932 36497 11966 36498
rect 12004 36497 12038 36498
rect 12076 36497 12110 36498
rect 12148 36497 12182 36498
rect 12220 36497 12254 36498
rect 12292 36497 12326 36498
rect 12364 36497 12398 36498
rect 12436 36497 12470 36498
rect 12508 36497 12542 36498
rect 12580 36497 12614 36498
rect 12652 36497 12686 36498
rect 12724 36497 12758 36498
rect 12796 36497 12830 36498
rect 12868 36497 12902 36498
rect 12940 36497 12974 36498
rect 13012 36497 13046 36498
rect 13084 36497 13118 36498
rect 13156 36497 13190 36498
rect 13228 36497 13262 36498
rect 13300 36497 13334 36498
rect 13372 36497 13406 36498
rect 13444 36497 13478 36498
rect 13516 36497 13550 36498
rect 13588 36497 13622 36498
rect 13660 36497 13694 36498
rect 13732 36497 13766 36498
rect 13804 36497 13838 36498
rect 13876 36497 13910 36498
rect 13948 36497 13982 36498
rect 14020 36497 14054 36498
rect 14092 36497 14126 36498
rect 14164 36497 14198 36498
rect 14236 36497 14270 36498
rect 14308 36497 14342 36498
rect 14380 36497 14414 36498
rect 556 36464 557 36497
rect 557 36464 590 36497
rect 628 36464 659 36497
rect 659 36464 662 36497
rect 700 36464 727 36497
rect 727 36464 734 36497
rect 772 36464 795 36497
rect 795 36464 806 36497
rect 844 36464 863 36497
rect 863 36464 878 36497
rect 916 36464 931 36497
rect 931 36464 950 36497
rect 988 36464 999 36497
rect 999 36464 1022 36497
rect 1060 36464 1067 36497
rect 1067 36464 1094 36497
rect 1132 36464 1135 36497
rect 1135 36464 1166 36497
rect 1204 36464 1237 36497
rect 1237 36464 1238 36497
rect 1276 36464 1305 36497
rect 1305 36464 1310 36497
rect 1348 36464 1373 36497
rect 1373 36464 1382 36497
rect 1420 36464 1441 36497
rect 1441 36464 1454 36497
rect 1492 36464 1509 36497
rect 1509 36464 1526 36497
rect 1564 36464 1577 36497
rect 1577 36464 1598 36497
rect 1636 36464 1645 36497
rect 1645 36464 1670 36497
rect 1708 36464 1713 36497
rect 1713 36464 1742 36497
rect 1780 36464 1781 36497
rect 1781 36464 1814 36497
rect 1852 36464 1883 36497
rect 1883 36464 1886 36497
rect 1924 36464 1951 36497
rect 1951 36464 1958 36497
rect 1996 36464 2019 36497
rect 2019 36464 2030 36497
rect 2068 36464 2087 36497
rect 2087 36464 2102 36497
rect 2140 36464 2155 36497
rect 2155 36464 2174 36497
rect 2212 36464 2223 36497
rect 2223 36464 2246 36497
rect 2284 36464 2291 36497
rect 2291 36464 2318 36497
rect 2356 36464 2359 36497
rect 2359 36464 2390 36497
rect 2428 36464 2461 36497
rect 2461 36464 2462 36497
rect 2500 36464 2529 36497
rect 2529 36464 2534 36497
rect 2572 36464 2597 36497
rect 2597 36464 2606 36497
rect 2644 36464 2665 36497
rect 2665 36464 2678 36497
rect 2716 36464 2733 36497
rect 2733 36464 2750 36497
rect 2788 36464 2801 36497
rect 2801 36464 2822 36497
rect 2860 36464 2869 36497
rect 2869 36464 2894 36497
rect 2932 36464 2937 36497
rect 2937 36464 2966 36497
rect 3004 36464 3005 36497
rect 3005 36464 3038 36497
rect 3076 36464 3107 36497
rect 3107 36464 3110 36497
rect 3148 36464 3175 36497
rect 3175 36464 3182 36497
rect 3220 36464 3243 36497
rect 3243 36464 3254 36497
rect 3292 36464 3311 36497
rect 3311 36464 3326 36497
rect 3364 36464 3379 36497
rect 3379 36464 3398 36497
rect 3436 36464 3447 36497
rect 3447 36464 3470 36497
rect 3508 36464 3515 36497
rect 3515 36464 3542 36497
rect 3580 36464 3583 36497
rect 3583 36464 3614 36497
rect 3652 36464 3685 36497
rect 3685 36464 3686 36497
rect 3724 36464 3753 36497
rect 3753 36464 3758 36497
rect 3796 36464 3821 36497
rect 3821 36464 3830 36497
rect 3868 36464 3889 36497
rect 3889 36464 3902 36497
rect 3940 36464 3957 36497
rect 3957 36464 3974 36497
rect 4012 36464 4025 36497
rect 4025 36464 4046 36497
rect 4084 36464 4093 36497
rect 4093 36464 4118 36497
rect 4156 36464 4161 36497
rect 4161 36464 4190 36497
rect 4228 36464 4229 36497
rect 4229 36464 4262 36497
rect 4300 36464 4331 36497
rect 4331 36464 4334 36497
rect 4372 36464 4399 36497
rect 4399 36464 4406 36497
rect 4444 36464 4467 36497
rect 4467 36464 4478 36497
rect 4516 36464 4535 36497
rect 4535 36464 4550 36497
rect 4588 36464 4603 36497
rect 4603 36464 4622 36497
rect 4660 36464 4671 36497
rect 4671 36464 4694 36497
rect 4732 36464 4739 36497
rect 4739 36464 4766 36497
rect 4804 36464 4807 36497
rect 4807 36464 4838 36497
rect 4876 36464 4909 36497
rect 4909 36464 4910 36497
rect 4948 36464 4977 36497
rect 4977 36464 4982 36497
rect 5020 36464 5045 36497
rect 5045 36464 5054 36497
rect 5092 36464 5113 36497
rect 5113 36464 5126 36497
rect 5164 36464 5181 36497
rect 5181 36464 5198 36497
rect 5236 36464 5249 36497
rect 5249 36464 5270 36497
rect 5308 36464 5317 36497
rect 5317 36464 5342 36497
rect 5380 36464 5385 36497
rect 5385 36464 5414 36497
rect 5452 36464 5453 36497
rect 5453 36464 5486 36497
rect 5524 36464 5555 36497
rect 5555 36464 5558 36497
rect 5596 36464 5623 36497
rect 5623 36464 5630 36497
rect 5668 36464 5691 36497
rect 5691 36464 5702 36497
rect 5740 36464 5759 36497
rect 5759 36464 5774 36497
rect 5812 36464 5827 36497
rect 5827 36464 5846 36497
rect 5884 36464 5895 36497
rect 5895 36464 5918 36497
rect 5956 36464 5963 36497
rect 5963 36464 5990 36497
rect 6028 36464 6031 36497
rect 6031 36464 6062 36497
rect 6100 36464 6133 36497
rect 6133 36464 6134 36497
rect 6172 36464 6201 36497
rect 6201 36464 6206 36497
rect 6244 36464 6269 36497
rect 6269 36464 6278 36497
rect 6316 36464 6337 36497
rect 6337 36464 6350 36497
rect 6388 36464 6405 36497
rect 6405 36464 6422 36497
rect 6460 36464 6473 36497
rect 6473 36464 6494 36497
rect 6532 36464 6541 36497
rect 6541 36464 6566 36497
rect 6604 36464 6609 36497
rect 6609 36464 6638 36497
rect 6676 36464 6677 36497
rect 6677 36464 6710 36497
rect 6748 36464 6779 36497
rect 6779 36464 6782 36497
rect 6820 36464 6847 36497
rect 6847 36464 6854 36497
rect 6892 36464 6915 36497
rect 6915 36464 6926 36497
rect 6964 36464 6983 36497
rect 6983 36464 6998 36497
rect 7036 36464 7051 36497
rect 7051 36464 7070 36497
rect 7108 36464 7119 36497
rect 7119 36464 7142 36497
rect 7180 36464 7187 36497
rect 7187 36464 7214 36497
rect 7252 36464 7255 36497
rect 7255 36464 7286 36497
rect 7324 36464 7357 36497
rect 7357 36464 7358 36497
rect 7396 36464 7425 36497
rect 7425 36464 7430 36497
rect 7468 36464 7493 36497
rect 7493 36464 7502 36497
rect 7540 36464 7561 36497
rect 7561 36464 7574 36497
rect 7612 36464 7629 36497
rect 7629 36464 7646 36497
rect 7684 36464 7697 36497
rect 7697 36464 7718 36497
rect 7756 36464 7765 36497
rect 7765 36464 7790 36497
rect 7828 36464 7833 36497
rect 7833 36464 7862 36497
rect 7900 36464 7901 36497
rect 7901 36464 7934 36497
rect 7972 36464 8003 36497
rect 8003 36464 8006 36497
rect 8044 36464 8071 36497
rect 8071 36464 8078 36497
rect 8116 36464 8139 36497
rect 8139 36464 8150 36497
rect 8188 36464 8207 36497
rect 8207 36464 8222 36497
rect 8260 36464 8275 36497
rect 8275 36464 8294 36497
rect 8332 36464 8343 36497
rect 8343 36464 8366 36497
rect 8404 36464 8411 36497
rect 8411 36464 8438 36497
rect 8476 36464 8479 36497
rect 8479 36464 8510 36497
rect 8548 36464 8581 36497
rect 8581 36464 8582 36497
rect 8620 36464 8649 36497
rect 8649 36464 8654 36497
rect 8692 36464 8717 36497
rect 8717 36464 8726 36497
rect 8764 36464 8785 36497
rect 8785 36464 8798 36497
rect 8836 36464 8853 36497
rect 8853 36464 8870 36497
rect 8908 36464 8921 36497
rect 8921 36464 8942 36497
rect 8980 36464 8989 36497
rect 8989 36464 9014 36497
rect 9052 36464 9057 36497
rect 9057 36464 9086 36497
rect 9124 36464 9125 36497
rect 9125 36464 9158 36497
rect 9196 36464 9227 36497
rect 9227 36464 9230 36497
rect 9268 36464 9295 36497
rect 9295 36464 9302 36497
rect 9340 36464 9363 36497
rect 9363 36464 9374 36497
rect 9412 36464 9431 36497
rect 9431 36464 9446 36497
rect 9484 36464 9499 36497
rect 9499 36464 9518 36497
rect 9556 36464 9567 36497
rect 9567 36464 9590 36497
rect 9628 36464 9635 36497
rect 9635 36464 9662 36497
rect 9700 36464 9703 36497
rect 9703 36464 9734 36497
rect 9772 36464 9805 36497
rect 9805 36464 9806 36497
rect 9844 36464 9873 36497
rect 9873 36464 9878 36497
rect 9916 36464 9941 36497
rect 9941 36464 9950 36497
rect 9988 36464 10009 36497
rect 10009 36464 10022 36497
rect 10060 36464 10077 36497
rect 10077 36464 10094 36497
rect 10132 36464 10145 36497
rect 10145 36464 10166 36497
rect 10204 36464 10213 36497
rect 10213 36464 10238 36497
rect 10276 36464 10281 36497
rect 10281 36464 10310 36497
rect 10348 36464 10349 36497
rect 10349 36464 10382 36497
rect 10420 36464 10451 36497
rect 10451 36464 10454 36497
rect 10492 36464 10519 36497
rect 10519 36464 10526 36497
rect 10564 36464 10587 36497
rect 10587 36464 10598 36497
rect 10636 36464 10655 36497
rect 10655 36464 10670 36497
rect 10708 36464 10723 36497
rect 10723 36464 10742 36497
rect 10780 36464 10791 36497
rect 10791 36464 10814 36497
rect 10852 36464 10859 36497
rect 10859 36464 10886 36497
rect 10924 36464 10927 36497
rect 10927 36464 10958 36497
rect 10996 36464 11029 36497
rect 11029 36464 11030 36497
rect 11068 36464 11097 36497
rect 11097 36464 11102 36497
rect 11140 36464 11165 36497
rect 11165 36464 11174 36497
rect 11212 36464 11233 36497
rect 11233 36464 11246 36497
rect 11284 36464 11301 36497
rect 11301 36464 11318 36497
rect 11356 36464 11369 36497
rect 11369 36464 11390 36497
rect 11428 36464 11437 36497
rect 11437 36464 11462 36497
rect 11500 36464 11505 36497
rect 11505 36464 11534 36497
rect 11572 36464 11573 36497
rect 11573 36464 11606 36497
rect 11644 36464 11675 36497
rect 11675 36464 11678 36497
rect 11716 36464 11743 36497
rect 11743 36464 11750 36497
rect 11788 36464 11811 36497
rect 11811 36464 11822 36497
rect 11860 36464 11879 36497
rect 11879 36464 11894 36497
rect 11932 36464 11947 36497
rect 11947 36464 11966 36497
rect 12004 36464 12015 36497
rect 12015 36464 12038 36497
rect 12076 36464 12083 36497
rect 12083 36464 12110 36497
rect 12148 36464 12151 36497
rect 12151 36464 12182 36497
rect 12220 36464 12253 36497
rect 12253 36464 12254 36497
rect 12292 36464 12321 36497
rect 12321 36464 12326 36497
rect 12364 36464 12389 36497
rect 12389 36464 12398 36497
rect 12436 36464 12457 36497
rect 12457 36464 12470 36497
rect 12508 36464 12525 36497
rect 12525 36464 12542 36497
rect 12580 36464 12593 36497
rect 12593 36464 12614 36497
rect 12652 36464 12661 36497
rect 12661 36464 12686 36497
rect 12724 36464 12729 36497
rect 12729 36464 12758 36497
rect 12796 36464 12797 36497
rect 12797 36464 12830 36497
rect 12868 36464 12899 36497
rect 12899 36464 12902 36497
rect 12940 36464 12967 36497
rect 12967 36464 12974 36497
rect 13012 36464 13035 36497
rect 13035 36464 13046 36497
rect 13084 36464 13103 36497
rect 13103 36464 13118 36497
rect 13156 36464 13171 36497
rect 13171 36464 13190 36497
rect 13228 36464 13239 36497
rect 13239 36464 13262 36497
rect 13300 36464 13307 36497
rect 13307 36464 13334 36497
rect 13372 36464 13375 36497
rect 13375 36464 13406 36497
rect 13444 36464 13477 36497
rect 13477 36464 13478 36497
rect 13516 36464 13545 36497
rect 13545 36464 13550 36497
rect 13588 36464 13613 36497
rect 13613 36464 13622 36497
rect 13660 36464 13681 36497
rect 13681 36464 13694 36497
rect 13732 36464 13749 36497
rect 13749 36464 13766 36497
rect 13804 36464 13817 36497
rect 13817 36464 13838 36497
rect 13876 36464 13885 36497
rect 13885 36464 13910 36497
rect 13948 36464 13953 36497
rect 13953 36464 13982 36497
rect 14020 36464 14021 36497
rect 14021 36464 14054 36497
rect 14092 36464 14123 36497
rect 14123 36464 14126 36497
rect 14164 36464 14191 36497
rect 14191 36464 14198 36497
rect 14236 36464 14259 36497
rect 14259 36464 14270 36497
rect 14308 36464 14327 36497
rect 14327 36464 14342 36497
rect 14380 36464 14395 36497
rect 14395 36464 14414 36497
rect 320 36428 354 36462
rect 14614 36427 14648 36461
rect 320 36254 346 36281
rect 346 36254 354 36281
rect 320 36247 354 36254
rect 320 36186 346 36209
rect 346 36186 354 36209
rect 320 36175 354 36186
rect 14614 36260 14641 36278
rect 14641 36260 14648 36278
rect 14614 36244 14648 36260
rect 320 36118 346 36137
rect 346 36118 354 36137
rect 320 36103 354 36118
rect 320 36050 346 36065
rect 346 36050 354 36065
rect 320 36031 354 36050
rect 320 35982 346 35993
rect 346 35982 354 35993
rect 320 35959 354 35982
rect 320 35914 346 35921
rect 346 35914 354 35921
rect 320 35887 354 35914
rect 320 35846 346 35849
rect 346 35846 354 35849
rect 320 35815 354 35846
rect 320 35744 354 35777
rect 320 35743 346 35744
rect 346 35743 354 35744
rect 320 35676 354 35705
rect 320 35671 346 35676
rect 346 35671 354 35676
rect 320 35608 354 35633
rect 320 35599 346 35608
rect 346 35599 354 35608
rect 320 35540 354 35561
rect 320 35527 346 35540
rect 346 35527 354 35540
rect 320 35472 354 35489
rect 320 35455 346 35472
rect 346 35455 354 35472
rect 320 35404 354 35417
rect 320 35383 346 35404
rect 346 35383 354 35404
rect 320 35336 354 35345
rect 320 35311 346 35336
rect 346 35311 354 35336
rect 320 35268 354 35273
rect 320 35239 346 35268
rect 346 35239 354 35268
rect 320 35200 354 35201
rect 320 35167 346 35200
rect 346 35167 354 35200
rect 320 35098 346 35129
rect 346 35098 354 35129
rect 320 35095 354 35098
rect 320 35030 346 35057
rect 346 35030 354 35057
rect 320 35023 354 35030
rect 320 34962 346 34985
rect 346 34962 354 34985
rect 320 34951 354 34962
rect 320 34894 346 34913
rect 346 34894 354 34913
rect 320 34879 354 34894
rect 320 34826 346 34841
rect 346 34826 354 34841
rect 320 34807 354 34826
rect 320 34758 346 34769
rect 346 34758 354 34769
rect 320 34735 354 34758
rect 320 34690 346 34697
rect 346 34690 354 34697
rect 320 34663 354 34690
rect 320 34622 346 34625
rect 346 34622 354 34625
rect 320 34591 354 34622
rect 320 34520 354 34553
rect 320 34519 346 34520
rect 346 34519 354 34520
rect 320 34452 354 34481
rect 320 34447 346 34452
rect 346 34447 354 34452
rect 320 34384 354 34409
rect 320 34375 346 34384
rect 346 34375 354 34384
rect 320 34316 354 34337
rect 320 34303 346 34316
rect 346 34303 354 34316
rect 320 34248 354 34265
rect 320 34231 346 34248
rect 346 34231 354 34248
rect 320 34180 354 34193
rect 320 34159 346 34180
rect 346 34159 354 34180
rect 320 34112 354 34121
rect 320 34087 346 34112
rect 346 34087 354 34112
rect 320 34044 354 34049
rect 320 34015 346 34044
rect 346 34015 354 34044
rect 320 33976 354 33977
rect 320 33943 346 33976
rect 346 33943 354 33976
rect 320 33874 346 33905
rect 346 33874 354 33905
rect 320 33871 354 33874
rect 320 33806 346 33833
rect 346 33806 354 33833
rect 320 33799 354 33806
rect 320 33738 346 33761
rect 346 33738 354 33761
rect 320 33727 354 33738
rect 320 33670 346 33689
rect 346 33670 354 33689
rect 320 33655 354 33670
rect 320 33602 346 33617
rect 346 33602 354 33617
rect 320 33583 354 33602
rect 320 33534 346 33545
rect 346 33534 354 33545
rect 320 33511 354 33534
rect 320 33466 346 33473
rect 346 33466 354 33473
rect 320 33439 354 33466
rect 320 33398 346 33401
rect 346 33398 354 33401
rect 320 33367 354 33398
rect 320 33296 354 33329
rect 320 33295 346 33296
rect 346 33295 354 33296
rect 320 33228 354 33257
rect 320 33223 346 33228
rect 346 33223 354 33228
rect 320 33160 354 33185
rect 320 33151 346 33160
rect 346 33151 354 33160
rect 320 33092 354 33113
rect 320 33079 346 33092
rect 346 33079 354 33092
rect 320 33024 354 33041
rect 320 33007 346 33024
rect 346 33007 354 33024
rect 320 32956 354 32969
rect 320 32935 346 32956
rect 346 32935 354 32956
rect 320 32888 354 32897
rect 320 32863 346 32888
rect 346 32863 354 32888
rect 320 32820 354 32825
rect 320 32791 346 32820
rect 346 32791 354 32820
rect 320 32752 354 32753
rect 320 32719 346 32752
rect 346 32719 354 32752
rect 320 32650 346 32681
rect 346 32650 354 32681
rect 320 32647 354 32650
rect 320 32582 346 32609
rect 346 32582 354 32609
rect 320 32575 354 32582
rect 320 32514 346 32537
rect 346 32514 354 32537
rect 320 32503 354 32514
rect 320 32446 346 32465
rect 346 32446 354 32465
rect 320 32431 354 32446
rect 320 32378 346 32393
rect 346 32378 354 32393
rect 320 32359 354 32378
rect 320 32310 346 32321
rect 346 32310 354 32321
rect 320 32287 354 32310
rect 320 32242 346 32249
rect 346 32242 354 32249
rect 320 32215 354 32242
rect 320 32174 346 32177
rect 346 32174 354 32177
rect 320 32143 354 32174
rect 320 32072 354 32105
rect 320 32071 346 32072
rect 346 32071 354 32072
rect 320 32004 354 32033
rect 320 31999 346 32004
rect 346 31999 354 32004
rect 320 31936 354 31961
rect 320 31927 346 31936
rect 346 31927 354 31936
rect 320 31868 354 31889
rect 320 31855 346 31868
rect 346 31855 354 31868
rect 320 31800 354 31817
rect 320 31783 346 31800
rect 346 31783 354 31800
rect 320 31732 354 31745
rect 320 31711 346 31732
rect 346 31711 354 31732
rect 320 31664 354 31673
rect 320 31639 346 31664
rect 346 31639 354 31664
rect 320 31596 354 31601
rect 320 31567 346 31596
rect 346 31567 354 31596
rect 320 31528 354 31529
rect 320 31495 346 31528
rect 346 31495 354 31528
rect 320 31426 346 31457
rect 346 31426 354 31457
rect 320 31423 354 31426
rect 320 31358 346 31385
rect 346 31358 354 31385
rect 320 31351 354 31358
rect 320 31290 346 31313
rect 346 31290 354 31313
rect 320 31279 354 31290
rect 320 31222 346 31241
rect 346 31222 354 31241
rect 320 31207 354 31222
rect 320 31154 346 31169
rect 346 31154 354 31169
rect 320 31135 354 31154
rect 320 31086 346 31097
rect 346 31086 354 31097
rect 320 31063 354 31086
rect 320 31018 346 31025
rect 346 31018 354 31025
rect 320 30991 354 31018
rect 320 30950 346 30953
rect 346 30950 354 30953
rect 320 30919 354 30950
rect 320 30848 354 30881
rect 320 30847 346 30848
rect 346 30847 354 30848
rect 320 30780 354 30809
rect 320 30775 346 30780
rect 346 30775 354 30780
rect 320 30712 354 30737
rect 320 30703 346 30712
rect 346 30703 354 30712
rect 320 30644 354 30665
rect 320 30631 346 30644
rect 346 30631 354 30644
rect 320 30576 354 30593
rect 320 30559 346 30576
rect 346 30559 354 30576
rect 320 30508 354 30521
rect 320 30487 346 30508
rect 346 30487 354 30508
rect 320 30440 354 30449
rect 320 30415 346 30440
rect 346 30415 354 30440
rect 320 30372 354 30377
rect 320 30343 346 30372
rect 346 30343 354 30372
rect 320 30304 354 30305
rect 320 30271 346 30304
rect 346 30271 354 30304
rect 320 30202 346 30233
rect 346 30202 354 30233
rect 320 30199 354 30202
rect 320 30134 346 30161
rect 346 30134 354 30161
rect 320 30127 354 30134
rect 320 30066 346 30089
rect 346 30066 354 30089
rect 320 30055 354 30066
rect 320 29998 346 30017
rect 346 29998 354 30017
rect 320 29983 354 29998
rect 320 29930 346 29945
rect 346 29930 354 29945
rect 320 29911 354 29930
rect 320 29862 346 29873
rect 346 29862 354 29873
rect 320 29839 354 29862
rect 320 29794 346 29801
rect 346 29794 354 29801
rect 320 29767 354 29794
rect 320 29726 346 29729
rect 346 29726 354 29729
rect 320 29695 354 29726
rect 320 29624 354 29657
rect 320 29623 346 29624
rect 346 29623 354 29624
rect 320 29556 354 29585
rect 320 29551 346 29556
rect 346 29551 354 29556
rect 320 29488 354 29513
rect 320 29479 346 29488
rect 346 29479 354 29488
rect 320 29420 354 29441
rect 320 29407 346 29420
rect 346 29407 354 29420
rect 320 29352 354 29369
rect 320 29335 346 29352
rect 346 29335 354 29352
rect 320 29284 354 29297
rect 320 29263 346 29284
rect 346 29263 354 29284
rect 320 29216 354 29225
rect 320 29191 346 29216
rect 346 29191 354 29216
rect 320 29148 354 29153
rect 320 29119 346 29148
rect 346 29119 354 29148
rect 320 29080 354 29081
rect 320 29047 346 29080
rect 346 29047 354 29080
rect 320 28978 346 29009
rect 346 28978 354 29009
rect 320 28975 354 28978
rect 320 28910 346 28937
rect 346 28910 354 28937
rect 320 28903 354 28910
rect 320 28842 346 28865
rect 346 28842 354 28865
rect 320 28831 354 28842
rect 320 28774 346 28793
rect 346 28774 354 28793
rect 320 28759 354 28774
rect 320 28706 346 28721
rect 346 28706 354 28721
rect 320 28687 354 28706
rect 320 28638 346 28649
rect 346 28638 354 28649
rect 320 28615 354 28638
rect 320 28570 346 28577
rect 346 28570 354 28577
rect 320 28543 354 28570
rect 320 28502 346 28505
rect 346 28502 354 28505
rect 320 28471 354 28502
rect 320 28400 354 28433
rect 320 28399 346 28400
rect 346 28399 354 28400
rect 320 28332 354 28361
rect 320 28327 346 28332
rect 346 28327 354 28332
rect 320 28264 354 28289
rect 320 28255 346 28264
rect 346 28255 354 28264
rect 320 28196 354 28217
rect 320 28183 346 28196
rect 346 28183 354 28196
rect 320 28128 354 28145
rect 320 28111 346 28128
rect 346 28111 354 28128
rect 320 28060 354 28073
rect 320 28039 346 28060
rect 346 28039 354 28060
rect 320 27992 354 28001
rect 320 27967 346 27992
rect 346 27967 354 27992
rect 320 27924 354 27929
rect 320 27895 346 27924
rect 346 27895 354 27924
rect 320 27856 354 27857
rect 320 27823 346 27856
rect 346 27823 354 27856
rect 320 27754 346 27785
rect 346 27754 354 27785
rect 320 27751 354 27754
rect 320 27686 346 27713
rect 346 27686 354 27713
rect 320 27679 354 27686
rect 320 27618 346 27641
rect 346 27618 354 27641
rect 320 27607 354 27618
rect 320 27550 346 27569
rect 346 27550 354 27569
rect 320 27535 354 27550
rect 320 27482 346 27497
rect 346 27482 354 27497
rect 320 27463 354 27482
rect 320 27414 346 27425
rect 346 27414 354 27425
rect 320 27391 354 27414
rect 320 27346 346 27353
rect 346 27346 354 27353
rect 320 27319 354 27346
rect 320 27278 346 27281
rect 346 27278 354 27281
rect 320 27247 354 27278
rect 320 27176 354 27209
rect 320 27175 346 27176
rect 346 27175 354 27176
rect 320 27108 354 27137
rect 320 27103 346 27108
rect 346 27103 354 27108
rect 320 27040 354 27065
rect 320 27031 346 27040
rect 346 27031 354 27040
rect 320 26972 354 26993
rect 320 26959 346 26972
rect 346 26959 354 26972
rect 320 26904 354 26921
rect 320 26887 346 26904
rect 346 26887 354 26904
rect 320 26836 354 26849
rect 320 26815 346 26836
rect 346 26815 354 26836
rect 320 26768 354 26777
rect 320 26743 346 26768
rect 346 26743 354 26768
rect 320 26700 354 26705
rect 320 26671 346 26700
rect 346 26671 354 26700
rect 320 26632 354 26633
rect 320 26599 346 26632
rect 346 26599 354 26632
rect 320 26530 346 26561
rect 346 26530 354 26561
rect 320 26527 354 26530
rect 320 26462 346 26489
rect 346 26462 354 26489
rect 320 26455 354 26462
rect 320 26394 346 26417
rect 346 26394 354 26417
rect 320 26383 354 26394
rect 320 26326 346 26345
rect 346 26326 354 26345
rect 320 26311 354 26326
rect 320 26258 346 26273
rect 346 26258 354 26273
rect 320 26239 354 26258
rect 320 26190 346 26201
rect 346 26190 354 26201
rect 320 26167 354 26190
rect 320 26122 346 26129
rect 346 26122 354 26129
rect 320 26095 354 26122
rect 320 26054 346 26057
rect 346 26054 354 26057
rect 320 26023 354 26054
rect 320 25952 354 25985
rect 320 25951 346 25952
rect 346 25951 354 25952
rect 320 25884 354 25913
rect 320 25879 346 25884
rect 346 25879 354 25884
rect 320 25816 354 25841
rect 320 25807 346 25816
rect 346 25807 354 25816
rect 320 25748 354 25769
rect 320 25735 346 25748
rect 346 25735 354 25748
rect 320 25680 354 25697
rect 320 25663 346 25680
rect 346 25663 354 25680
rect 320 25612 354 25625
rect 320 25591 346 25612
rect 346 25591 354 25612
rect 320 25544 354 25553
rect 320 25519 346 25544
rect 346 25519 354 25544
rect 320 25476 354 25481
rect 320 25447 346 25476
rect 346 25447 354 25476
rect 320 25408 354 25409
rect 320 25375 346 25408
rect 346 25375 354 25408
rect 320 25306 346 25337
rect 346 25306 354 25337
rect 320 25303 354 25306
rect 320 25238 346 25265
rect 346 25238 354 25265
rect 320 25231 354 25238
rect 320 25170 346 25193
rect 346 25170 354 25193
rect 320 25159 354 25170
rect 320 25102 346 25121
rect 346 25102 354 25121
rect 320 25087 354 25102
rect 320 25034 346 25049
rect 346 25034 354 25049
rect 320 25015 354 25034
rect 320 24966 346 24977
rect 346 24966 354 24977
rect 320 24943 354 24966
rect 320 24898 346 24905
rect 346 24898 354 24905
rect 320 24871 354 24898
rect 320 24830 346 24833
rect 346 24830 354 24833
rect 320 24799 354 24830
rect 320 24728 354 24761
rect 320 24727 346 24728
rect 346 24727 354 24728
rect 320 24660 354 24689
rect 320 24655 346 24660
rect 346 24655 354 24660
rect 320 24592 354 24617
rect 320 24583 346 24592
rect 346 24583 354 24592
rect 320 24524 354 24545
rect 320 24511 346 24524
rect 346 24511 354 24524
rect 320 24456 354 24473
rect 320 24439 346 24456
rect 346 24439 354 24456
rect 320 24388 354 24401
rect 320 24367 346 24388
rect 346 24367 354 24388
rect 320 24320 354 24329
rect 320 24295 346 24320
rect 346 24295 354 24320
rect 320 24252 354 24257
rect 320 24223 346 24252
rect 346 24223 354 24252
rect 320 24184 354 24185
rect 320 24151 346 24184
rect 346 24151 354 24184
rect 320 24082 346 24113
rect 346 24082 354 24113
rect 320 24079 354 24082
rect 320 24014 346 24041
rect 346 24014 354 24041
rect 320 24007 354 24014
rect 320 23946 346 23969
rect 346 23946 354 23969
rect 320 23935 354 23946
rect 320 23878 346 23897
rect 346 23878 354 23897
rect 320 23863 354 23878
rect 320 23810 346 23825
rect 346 23810 354 23825
rect 320 23791 354 23810
rect 320 23742 346 23753
rect 346 23742 354 23753
rect 320 23719 354 23742
rect 320 23674 346 23681
rect 346 23674 354 23681
rect 320 23647 354 23674
rect 320 23606 346 23609
rect 346 23606 354 23609
rect 320 23575 354 23606
rect 320 23504 354 23537
rect 320 23503 346 23504
rect 346 23503 354 23504
rect 320 23436 354 23465
rect 320 23431 346 23436
rect 346 23431 354 23436
rect 320 23368 354 23393
rect 320 23359 346 23368
rect 346 23359 354 23368
rect 320 23300 354 23321
rect 320 23287 346 23300
rect 346 23287 354 23300
rect 320 23232 354 23249
rect 320 23215 346 23232
rect 346 23215 354 23232
rect 320 23164 354 23177
rect 320 23143 346 23164
rect 346 23143 354 23164
rect 320 23096 354 23105
rect 320 23071 346 23096
rect 346 23071 354 23096
rect 320 23028 354 23033
rect 320 22999 346 23028
rect 346 22999 354 23028
rect 320 22960 354 22961
rect 320 22927 346 22960
rect 346 22927 354 22960
rect 320 22858 346 22889
rect 346 22858 354 22889
rect 320 22855 354 22858
rect 320 22790 346 22817
rect 346 22790 354 22817
rect 320 22783 354 22790
rect 320 22722 346 22745
rect 346 22722 354 22745
rect 320 22711 354 22722
rect 320 22654 346 22673
rect 346 22654 354 22673
rect 320 22639 354 22654
rect 320 22586 346 22601
rect 346 22586 354 22601
rect 320 22567 354 22586
rect 320 22518 346 22529
rect 346 22518 354 22529
rect 320 22495 354 22518
rect 320 22450 346 22457
rect 346 22450 354 22457
rect 320 22423 354 22450
rect 320 22382 346 22385
rect 346 22382 354 22385
rect 320 22351 354 22382
rect 320 22280 354 22313
rect 320 22279 346 22280
rect 346 22279 354 22280
rect 320 22212 354 22241
rect 320 22207 346 22212
rect 346 22207 354 22212
rect 320 22144 354 22169
rect 320 22135 346 22144
rect 346 22135 354 22144
rect 320 22076 354 22097
rect 320 22063 346 22076
rect 346 22063 354 22076
rect 320 22008 354 22025
rect 320 21991 346 22008
rect 346 21991 354 22008
rect 320 21940 354 21953
rect 320 21919 346 21940
rect 346 21919 354 21940
rect 320 21872 354 21881
rect 320 21847 346 21872
rect 346 21847 354 21872
rect 320 21804 354 21809
rect 320 21775 346 21804
rect 346 21775 354 21804
rect 320 21736 354 21737
rect 320 21703 346 21736
rect 346 21703 354 21736
rect 320 21634 346 21665
rect 346 21634 354 21665
rect 320 21631 354 21634
rect 320 21566 346 21593
rect 346 21566 354 21593
rect 320 21559 354 21566
rect 320 21498 346 21521
rect 346 21498 354 21521
rect 320 21487 354 21498
rect 320 21430 346 21449
rect 346 21430 354 21449
rect 320 21415 354 21430
rect 320 21362 346 21377
rect 346 21362 354 21377
rect 320 21343 354 21362
rect 320 21294 346 21305
rect 346 21294 354 21305
rect 320 21271 354 21294
rect 320 21226 346 21233
rect 346 21226 354 21233
rect 320 21199 354 21226
rect 320 21158 346 21161
rect 346 21158 354 21161
rect 320 21127 354 21158
rect 320 21056 354 21089
rect 320 21055 346 21056
rect 346 21055 354 21056
rect 320 20988 354 21017
rect 320 20983 346 20988
rect 346 20983 354 20988
rect 320 20920 354 20945
rect 320 20911 346 20920
rect 346 20911 354 20920
rect 320 20852 354 20873
rect 320 20839 346 20852
rect 346 20839 354 20852
rect 320 20784 354 20801
rect 320 20767 346 20784
rect 346 20767 354 20784
rect 320 20716 354 20729
rect 320 20695 346 20716
rect 346 20695 354 20716
rect 320 20648 354 20657
rect 320 20623 346 20648
rect 346 20623 354 20648
rect 320 20580 354 20585
rect 320 20551 346 20580
rect 346 20551 354 20580
rect 320 20512 354 20513
rect 320 20479 346 20512
rect 346 20479 354 20512
rect 320 20410 346 20441
rect 346 20410 354 20441
rect 320 20407 354 20410
rect 320 20342 346 20369
rect 346 20342 354 20369
rect 320 20335 354 20342
rect 320 20274 346 20297
rect 346 20274 354 20297
rect 320 20263 354 20274
rect 320 20206 346 20225
rect 346 20206 354 20225
rect 320 20191 354 20206
rect 320 20138 346 20153
rect 346 20138 354 20153
rect 320 20119 354 20138
rect 320 20070 346 20081
rect 346 20070 354 20081
rect 320 20047 354 20070
rect 320 20002 346 20009
rect 346 20002 354 20009
rect 320 19975 354 20002
rect 320 19934 346 19937
rect 346 19934 354 19937
rect 320 19903 354 19934
rect 320 19832 354 19865
rect 320 19831 346 19832
rect 346 19831 354 19832
rect 320 19764 354 19793
rect 320 19759 346 19764
rect 346 19759 354 19764
rect 320 19696 354 19721
rect 320 19687 346 19696
rect 346 19687 354 19696
rect 320 19628 354 19649
rect 320 19615 346 19628
rect 346 19615 354 19628
rect 320 19560 354 19577
rect 320 19543 346 19560
rect 346 19543 354 19560
rect 320 19492 354 19505
rect 320 19471 346 19492
rect 346 19471 354 19492
rect 320 19424 354 19433
rect 320 19399 346 19424
rect 346 19399 354 19424
rect 320 19356 354 19361
rect 320 19327 346 19356
rect 346 19327 354 19356
rect 320 19288 354 19289
rect 320 19255 346 19288
rect 346 19255 354 19288
rect 320 19186 346 19217
rect 346 19186 354 19217
rect 320 19183 354 19186
rect 320 19118 346 19145
rect 346 19118 354 19145
rect 320 19111 354 19118
rect 320 19050 346 19073
rect 346 19050 354 19073
rect 320 19039 354 19050
rect 320 18982 346 19001
rect 346 18982 354 19001
rect 320 18967 354 18982
rect 320 18914 346 18929
rect 346 18914 354 18929
rect 320 18895 354 18914
rect 320 18846 346 18857
rect 346 18846 354 18857
rect 320 18823 354 18846
rect 320 18778 346 18785
rect 346 18778 354 18785
rect 320 18751 354 18778
rect 320 18710 346 18713
rect 346 18710 354 18713
rect 320 18679 354 18710
rect 320 18608 354 18641
rect 320 18607 346 18608
rect 346 18607 354 18608
rect 320 18540 354 18569
rect 320 18535 346 18540
rect 346 18535 354 18540
rect 320 18472 354 18497
rect 320 18463 346 18472
rect 346 18463 354 18472
rect 320 18404 354 18425
rect 320 18391 346 18404
rect 346 18391 354 18404
rect 320 18336 354 18353
rect 320 18319 346 18336
rect 346 18319 354 18336
rect 320 18268 354 18281
rect 320 18247 346 18268
rect 346 18247 354 18268
rect 320 18200 354 18209
rect 320 18175 346 18200
rect 346 18175 354 18200
rect 320 18132 354 18137
rect 320 18103 346 18132
rect 346 18103 354 18132
rect 320 18064 354 18065
rect 320 18031 346 18064
rect 346 18031 354 18064
rect 320 17962 346 17993
rect 346 17962 354 17993
rect 320 17959 354 17962
rect 320 17894 346 17921
rect 346 17894 354 17921
rect 320 17887 354 17894
rect 320 17826 346 17849
rect 346 17826 354 17849
rect 320 17815 354 17826
rect 320 17758 346 17777
rect 346 17758 354 17777
rect 320 17743 354 17758
rect 320 17690 346 17705
rect 346 17690 354 17705
rect 320 17671 354 17690
rect 320 17622 346 17633
rect 346 17622 354 17633
rect 320 17599 354 17622
rect 320 17554 346 17561
rect 346 17554 354 17561
rect 320 17527 354 17554
rect 320 17486 346 17489
rect 346 17486 354 17489
rect 320 17455 354 17486
rect 320 17384 354 17417
rect 320 17383 346 17384
rect 346 17383 354 17384
rect 320 17316 354 17345
rect 320 17311 346 17316
rect 346 17311 354 17316
rect 320 17248 354 17273
rect 320 17239 346 17248
rect 346 17239 354 17248
rect 320 17180 354 17201
rect 320 17167 346 17180
rect 346 17167 354 17180
rect 320 17112 354 17129
rect 320 17095 346 17112
rect 346 17095 354 17112
rect 320 17044 354 17057
rect 320 17023 346 17044
rect 346 17023 354 17044
rect 320 16976 354 16985
rect 320 16951 346 16976
rect 346 16951 354 16976
rect 320 16908 354 16913
rect 320 16879 346 16908
rect 346 16879 354 16908
rect 320 16840 354 16841
rect 320 16807 346 16840
rect 346 16807 354 16840
rect 320 16738 346 16769
rect 346 16738 354 16769
rect 320 16735 354 16738
rect 320 16670 346 16697
rect 346 16670 354 16697
rect 320 16663 354 16670
rect 320 16602 346 16625
rect 346 16602 354 16625
rect 320 16591 354 16602
rect 320 16534 346 16553
rect 346 16534 354 16553
rect 320 16519 354 16534
rect 320 16466 346 16481
rect 346 16466 354 16481
rect 320 16447 354 16466
rect 320 16398 346 16409
rect 346 16398 354 16409
rect 320 16375 354 16398
rect 320 16330 346 16337
rect 346 16330 354 16337
rect 320 16303 354 16330
rect 320 16262 346 16265
rect 346 16262 354 16265
rect 320 16231 354 16262
rect 320 16160 354 16193
rect 320 16159 346 16160
rect 346 16159 354 16160
rect 320 16092 354 16121
rect 320 16087 346 16092
rect 346 16087 354 16092
rect 320 16024 354 16049
rect 320 16015 346 16024
rect 346 16015 354 16024
rect 320 15956 354 15977
rect 320 15943 346 15956
rect 346 15943 354 15956
rect 320 15888 354 15905
rect 320 15871 346 15888
rect 346 15871 354 15888
rect 320 15820 354 15833
rect 320 15799 346 15820
rect 346 15799 354 15820
rect 320 15752 354 15761
rect 320 15727 346 15752
rect 346 15727 354 15752
rect 320 15684 354 15689
rect 320 15655 346 15684
rect 346 15655 354 15684
rect 320 15616 354 15617
rect 320 15583 346 15616
rect 346 15583 354 15616
rect 320 15514 346 15545
rect 346 15514 354 15545
rect 320 15511 354 15514
rect 320 15446 346 15473
rect 346 15446 354 15473
rect 320 15439 354 15446
rect 320 15378 346 15401
rect 346 15378 354 15401
rect 320 15367 354 15378
rect 320 15310 346 15329
rect 346 15310 354 15329
rect 320 15295 354 15310
rect 320 15242 346 15257
rect 346 15242 354 15257
rect 320 15223 354 15242
rect 320 15174 346 15185
rect 346 15174 354 15185
rect 320 15151 354 15174
rect 320 15106 346 15113
rect 346 15106 354 15113
rect 320 15079 354 15106
rect 320 15038 346 15041
rect 346 15038 354 15041
rect 320 15007 354 15038
rect 320 14936 354 14969
rect 320 14935 346 14936
rect 346 14935 354 14936
rect 320 14868 354 14897
rect 320 14863 346 14868
rect 346 14863 354 14868
rect 320 14800 354 14825
rect 320 14791 346 14800
rect 346 14791 354 14800
rect 320 14732 354 14753
rect 320 14719 346 14732
rect 346 14719 354 14732
rect 1009 35969 1043 36003
rect 1081 35969 1115 36003
rect 1153 35969 1187 36003
rect 1225 35969 1259 36003
rect 1297 35969 1331 36003
rect 1369 35969 1403 36003
rect 1441 35969 1475 36003
rect 1513 35969 1547 36003
rect 1585 35969 1619 36003
rect 1657 35969 1691 36003
rect 1729 35969 1763 36003
rect 1801 35969 1835 36003
rect 1873 35969 1907 36003
rect 1945 35969 1979 36003
rect 2017 35969 2051 36003
rect 2089 35969 2123 36003
rect 2161 35969 2195 36003
rect 2233 35969 2267 36003
rect 2305 35969 2339 36003
rect 2377 35969 2411 36003
rect 2449 35969 2483 36003
rect 2521 35969 2555 36003
rect 2593 35969 2627 36003
rect 2665 35969 2699 36003
rect 2737 35969 2771 36003
rect 2809 35969 2843 36003
rect 2881 35969 2915 36003
rect 2953 35969 2987 36003
rect 3025 35969 3059 36003
rect 3097 35969 3131 36003
rect 3169 35969 3203 36003
rect 3241 35969 3275 36003
rect 3313 35969 3347 36003
rect 3385 35969 3419 36003
rect 3457 35969 3491 36003
rect 3529 35969 3563 36003
rect 3601 35969 3635 36003
rect 3673 35969 3707 36003
rect 3745 35969 3779 36003
rect 3817 35969 3851 36003
rect 3889 35969 3923 36003
rect 3961 35969 3995 36003
rect 4033 35969 4067 36003
rect 4105 35969 4139 36003
rect 4177 35969 4211 36003
rect 4249 35969 4283 36003
rect 4321 35969 4355 36003
rect 4393 35969 4427 36003
rect 4465 35969 4499 36003
rect 4537 35969 4571 36003
rect 4609 35969 4643 36003
rect 4681 35969 4715 36003
rect 4753 35969 4787 36003
rect 4825 35969 4859 36003
rect 4897 35969 4931 36003
rect 4969 35969 5003 36003
rect 5041 35969 5075 36003
rect 5113 35969 5147 36003
rect 5185 35969 5219 36003
rect 5257 35969 5291 36003
rect 5329 35969 5363 36003
rect 5401 35969 5435 36003
rect 5473 35969 5507 36003
rect 5545 35969 5579 36003
rect 5617 35969 5651 36003
rect 5689 35969 5723 36003
rect 5761 35969 5795 36003
rect 5833 35969 5867 36003
rect 5905 35969 5939 36003
rect 5977 35969 6011 36003
rect 6049 35969 6083 36003
rect 6121 35969 6155 36003
rect 6193 35969 6227 36003
rect 6265 35969 6299 36003
rect 6337 35969 6371 36003
rect 6409 35969 6443 36003
rect 6481 35969 6515 36003
rect 6553 35969 6587 36003
rect 6625 35969 6659 36003
rect 6697 35969 6731 36003
rect 6769 35969 6803 36003
rect 6841 35969 6875 36003
rect 6913 35969 6947 36003
rect 6985 35969 7019 36003
rect 7057 35969 7091 36003
rect 7129 35969 7163 36003
rect 7201 35969 7235 36003
rect 7273 35969 7307 36003
rect 7345 35969 7379 36003
rect 7417 35969 7451 36003
rect 7489 35969 7523 36003
rect 7561 35969 7595 36003
rect 7633 35969 7667 36003
rect 7705 35969 7739 36003
rect 7777 35969 7811 36003
rect 7849 35969 7883 36003
rect 7921 35969 7955 36003
rect 7993 35969 8027 36003
rect 8065 35969 8099 36003
rect 8137 35969 8171 36003
rect 8209 35969 8243 36003
rect 8281 35969 8315 36003
rect 8353 35969 8387 36003
rect 8425 35969 8459 36003
rect 8497 35969 8531 36003
rect 8569 35969 8603 36003
rect 8641 35969 8675 36003
rect 8713 35969 8747 36003
rect 8785 35969 8819 36003
rect 8857 35969 8891 36003
rect 8929 35969 8963 36003
rect 9001 35969 9035 36003
rect 9073 35969 9107 36003
rect 9145 35969 9179 36003
rect 9217 35969 9251 36003
rect 9289 35969 9323 36003
rect 9361 35969 9395 36003
rect 9433 35969 9467 36003
rect 9505 35969 9539 36003
rect 9577 35969 9611 36003
rect 9649 35969 9683 36003
rect 9721 35969 9755 36003
rect 9793 35969 9827 36003
rect 9865 35969 9899 36003
rect 9937 35969 9971 36003
rect 10009 35969 10043 36003
rect 10081 35969 10115 36003
rect 10153 35969 10187 36003
rect 10225 35969 10259 36003
rect 10297 35969 10331 36003
rect 10369 35969 10403 36003
rect 10441 35969 10475 36003
rect 10513 35969 10547 36003
rect 10585 35969 10619 36003
rect 10657 35969 10691 36003
rect 10729 35969 10763 36003
rect 10801 35969 10835 36003
rect 10873 35969 10907 36003
rect 10945 35969 10979 36003
rect 11017 35969 11051 36003
rect 11089 35969 11123 36003
rect 11161 35969 11195 36003
rect 11233 35969 11267 36003
rect 11305 35969 11339 36003
rect 11377 35969 11411 36003
rect 11449 35969 11483 36003
rect 11521 35969 11555 36003
rect 11593 35969 11627 36003
rect 11665 35969 11699 36003
rect 11737 35969 11771 36003
rect 11809 35969 11843 36003
rect 11881 35969 11915 36003
rect 11953 35969 11987 36003
rect 12025 35969 12059 36003
rect 12097 35969 12131 36003
rect 12169 35969 12203 36003
rect 12241 35969 12275 36003
rect 12313 35969 12347 36003
rect 12385 35969 12419 36003
rect 12457 35969 12491 36003
rect 12529 35969 12563 36003
rect 12601 35969 12635 36003
rect 12673 35969 12707 36003
rect 12745 35969 12779 36003
rect 12817 35969 12851 36003
rect 12889 35969 12923 36003
rect 12961 35969 12995 36003
rect 13033 35969 13067 36003
rect 13105 35969 13139 36003
rect 13177 35969 13211 36003
rect 13249 35969 13283 36003
rect 13321 35969 13355 36003
rect 13393 35969 13427 36003
rect 13465 35969 13499 36003
rect 13537 35969 13571 36003
rect 13609 35969 13643 36003
rect 13681 35969 13715 36003
rect 13753 35969 13787 36003
rect 13825 35969 13859 36003
rect 13897 35969 13931 36003
rect 13969 35969 14003 36003
rect 807 35866 841 35900
rect 807 35794 841 35828
rect 14122 35787 14156 35821
rect 807 35722 841 35756
rect 14122 35715 14156 35749
rect 807 35650 841 35684
rect 14122 35643 14156 35677
rect 807 35578 841 35612
rect 14122 35571 14156 35605
rect 807 35506 841 35540
rect 14122 35499 14156 35533
rect 807 35434 841 35468
rect 14122 35427 14156 35461
rect 807 35362 841 35396
rect 14122 35355 14156 35389
rect 807 35290 841 35324
rect 14122 35283 14156 35317
rect 807 35218 841 35252
rect 14122 35211 14156 35245
rect 807 35146 841 35180
rect 14122 35139 14156 35173
rect 807 35074 841 35108
rect 14122 35067 14156 35101
rect 807 35002 841 35036
rect 14122 34995 14156 35029
rect 807 34930 841 34964
rect 14122 34923 14156 34957
rect 807 34858 841 34892
rect 14122 34851 14156 34885
rect 807 34786 841 34820
rect 807 34714 841 34748
rect 14122 34779 14156 34813
rect 807 34642 841 34676
rect 807 34570 841 34604
rect 807 34498 841 34532
rect 807 34426 841 34460
rect 807 34354 841 34388
rect 807 34282 841 34316
rect 807 34210 841 34244
rect 807 34138 841 34172
rect 807 34066 841 34100
rect 807 33994 841 34028
rect 807 33922 841 33956
rect 807 33850 841 33884
rect 807 33778 841 33812
rect 807 33706 841 33740
rect 807 33634 841 33668
rect 807 33562 841 33596
rect 807 33490 841 33524
rect 807 33418 841 33452
rect 807 33346 841 33380
rect 807 33274 841 33308
rect 807 33202 841 33236
rect 807 33130 841 33164
rect 807 33058 841 33092
rect 807 32986 841 33020
rect 807 32914 841 32948
rect 807 32842 841 32876
rect 807 32770 841 32804
rect 807 32698 841 32732
rect 807 32626 841 32660
rect 807 32554 841 32588
rect 807 32482 841 32516
rect 807 32410 841 32444
rect 807 32338 841 32372
rect 807 32266 841 32300
rect 807 32194 841 32228
rect 807 32122 841 32156
rect 807 32050 841 32084
rect 807 31978 841 32012
rect 807 31906 841 31940
rect 807 31834 841 31868
rect 807 31762 841 31796
rect 807 31690 841 31724
rect 807 31618 841 31652
rect 807 31546 841 31580
rect 807 31474 841 31508
rect 807 31402 841 31436
rect 807 31330 841 31364
rect 807 31258 841 31292
rect 807 31186 841 31220
rect 807 31114 841 31148
rect 807 31042 841 31076
rect 807 30970 841 31004
rect 807 30898 841 30932
rect 807 30826 841 30860
rect 807 30754 841 30788
rect 807 30682 841 30716
rect 807 30610 841 30644
rect 807 30538 841 30572
rect 807 30466 841 30500
rect 807 30394 841 30428
rect 807 30322 841 30356
rect 807 30250 841 30284
rect 807 30178 841 30212
rect 807 30106 841 30140
rect 807 30034 841 30068
rect 807 29962 841 29996
rect 807 29890 841 29924
rect 807 29818 841 29852
rect 807 29746 841 29780
rect 807 29674 841 29708
rect 807 29602 841 29636
rect 807 29530 841 29564
rect 807 29458 841 29492
rect 807 29386 841 29420
rect 807 29314 841 29348
rect 807 29242 841 29276
rect 807 29170 841 29204
rect 807 29098 841 29132
rect 807 29026 841 29060
rect 807 28954 841 28988
rect 807 28882 841 28916
rect 807 28810 841 28844
rect 807 28738 841 28772
rect 807 28666 841 28700
rect 807 28594 841 28628
rect 807 28522 841 28556
rect 807 28450 841 28484
rect 807 28378 841 28412
rect 807 28306 841 28340
rect 807 28234 841 28268
rect 807 28162 841 28196
rect 807 28090 841 28124
rect 807 28018 841 28052
rect 807 27946 841 27980
rect 807 27874 841 27908
rect 807 27802 841 27836
rect 807 27730 841 27764
rect 807 27658 841 27692
rect 807 27586 841 27620
rect 807 27514 841 27548
rect 807 27442 841 27476
rect 807 27370 841 27404
rect 807 27298 841 27332
rect 807 27226 841 27260
rect 807 27154 841 27188
rect 807 27082 841 27116
rect 807 27010 841 27044
rect 807 26938 841 26972
rect 807 26866 841 26900
rect 807 26794 841 26828
rect 807 26722 841 26756
rect 807 26650 841 26684
rect 807 26578 841 26612
rect 807 26506 841 26540
rect 807 26434 841 26468
rect 807 26362 841 26396
rect 807 26290 841 26324
rect 807 26218 841 26252
rect 807 26146 841 26180
rect 807 26074 841 26108
rect 807 26002 841 26036
rect 807 25930 841 25964
rect 807 25858 841 25892
rect 807 25786 841 25820
rect 807 25714 841 25748
rect 807 25642 841 25676
rect 807 25570 841 25604
rect 807 25498 841 25532
rect 807 25426 841 25460
rect 807 25354 841 25388
rect 807 25282 841 25316
rect 807 25210 841 25244
rect 807 25138 841 25172
rect 807 25066 841 25100
rect 807 24994 841 25028
rect 807 24922 841 24956
rect 807 24850 841 24884
rect 807 24778 841 24812
rect 807 24706 841 24740
rect 807 24634 841 24668
rect 807 24562 841 24596
rect 807 24490 841 24524
rect 807 24418 841 24452
rect 807 24346 841 24380
rect 807 24274 841 24308
rect 807 24202 841 24236
rect 807 24130 841 24164
rect 807 24058 841 24092
rect 807 23986 841 24020
rect 807 23914 841 23948
rect 807 23842 841 23876
rect 807 23770 841 23804
rect 807 23698 841 23732
rect 807 23626 841 23660
rect 807 23554 841 23588
rect 807 23482 841 23516
rect 807 23410 841 23444
rect 807 23338 841 23372
rect 807 23266 841 23300
rect 807 23194 841 23228
rect 807 23122 841 23156
rect 807 23050 841 23084
rect 807 22978 841 23012
rect 807 22906 841 22940
rect 807 22834 841 22868
rect 807 22762 841 22796
rect 807 22690 841 22724
rect 807 22618 841 22652
rect 807 22546 841 22580
rect 807 22474 841 22508
rect 807 22402 841 22436
rect 807 22330 841 22364
rect 807 22258 841 22292
rect 807 22186 841 22220
rect 807 22114 841 22148
rect 807 22042 841 22076
rect 807 21970 841 22004
rect 807 21898 841 21932
rect 807 21826 841 21860
rect 807 21754 841 21788
rect 807 21682 841 21716
rect 807 21610 841 21644
rect 807 21538 841 21572
rect 807 21466 841 21500
rect 807 21394 841 21428
rect 807 21322 841 21356
rect 807 21250 841 21284
rect 807 21178 841 21212
rect 807 21106 841 21140
rect 807 21034 841 21068
rect 807 20962 841 20996
rect 807 20890 841 20924
rect 807 20818 841 20852
rect 807 20746 841 20780
rect 807 20674 841 20708
rect 807 20602 841 20636
rect 807 20530 841 20564
rect 807 20458 841 20492
rect 807 20386 841 20420
rect 807 20314 841 20348
rect 807 20242 841 20276
rect 807 20170 841 20204
rect 807 20098 841 20132
rect 807 20026 841 20060
rect 807 19954 841 19988
rect 807 19882 841 19916
rect 807 19810 841 19844
rect 807 19738 841 19772
rect 807 19666 841 19700
rect 807 19594 841 19628
rect 807 19522 841 19556
rect 807 19450 841 19484
rect 807 19378 841 19412
rect 807 19306 841 19340
rect 807 19234 841 19268
rect 807 19162 841 19196
rect 807 19090 841 19124
rect 807 19018 841 19052
rect 807 18946 841 18980
rect 807 18874 841 18908
rect 807 18802 841 18836
rect 807 18730 841 18764
rect 807 18658 841 18692
rect 807 18586 841 18620
rect 807 18514 841 18548
rect 807 18442 841 18476
rect 807 18370 841 18404
rect 807 18298 841 18332
rect 807 18226 841 18260
rect 807 18154 841 18188
rect 807 18082 841 18116
rect 807 18010 841 18044
rect 807 17938 841 17972
rect 807 17866 841 17900
rect 807 17794 841 17828
rect 807 17722 841 17756
rect 807 17650 841 17684
rect 807 17578 841 17612
rect 807 17506 841 17540
rect 807 17434 841 17468
rect 807 17362 841 17396
rect 807 17290 841 17324
rect 807 17218 841 17252
rect 807 17146 841 17180
rect 807 17074 841 17108
rect 807 17002 841 17036
rect 807 16930 841 16964
rect 807 16858 841 16892
rect 807 16786 841 16820
rect 807 16714 841 16748
rect 807 16642 841 16676
rect 807 16570 841 16604
rect 807 16498 841 16532
rect 807 16426 841 16460
rect 807 16354 841 16388
rect 807 16282 841 16316
rect 807 16210 841 16244
rect 807 16138 841 16172
rect 807 16066 841 16100
rect 807 15994 841 16028
rect 807 15922 841 15956
rect 807 15850 841 15884
rect 807 15778 841 15812
rect 807 15706 841 15740
rect 807 15634 841 15668
rect 807 15562 841 15596
rect 807 15490 841 15524
rect 807 15418 841 15452
rect 807 15346 841 15380
rect 807 15274 841 15308
rect 807 15202 841 15236
rect 1301 34645 1305 34679
rect 1305 34645 1335 34679
rect 1373 34645 1407 34679
rect 1445 34645 1475 34679
rect 1475 34645 1479 34679
rect 1517 34645 1543 34679
rect 1543 34645 1551 34679
rect 1589 34645 1611 34679
rect 1611 34645 1623 34679
rect 1661 34645 1679 34679
rect 1679 34645 1695 34679
rect 1733 34645 1747 34679
rect 1747 34645 1767 34679
rect 1805 34645 1815 34679
rect 1815 34645 1839 34679
rect 1877 34645 1883 34679
rect 1883 34645 1911 34679
rect 1949 34645 1951 34679
rect 1951 34645 1983 34679
rect 2021 34645 2053 34679
rect 2053 34645 2055 34679
rect 2093 34645 2121 34679
rect 2121 34645 2127 34679
rect 2165 34645 2189 34679
rect 2189 34645 2199 34679
rect 2237 34645 2257 34679
rect 2257 34645 2271 34679
rect 2309 34645 2325 34679
rect 2325 34645 2343 34679
rect 2381 34645 2393 34679
rect 2393 34645 2415 34679
rect 2453 34645 2461 34679
rect 2461 34645 2487 34679
rect 2525 34645 2529 34679
rect 2529 34645 2559 34679
rect 2597 34645 2631 34679
rect 2669 34645 2699 34679
rect 2699 34645 2703 34679
rect 2741 34645 2767 34679
rect 2767 34645 2775 34679
rect 2813 34645 2835 34679
rect 2835 34645 2847 34679
rect 2885 34645 2903 34679
rect 2903 34645 2919 34679
rect 2957 34645 2971 34679
rect 2971 34645 2991 34679
rect 3029 34645 3039 34679
rect 3039 34645 3063 34679
rect 3101 34645 3107 34679
rect 3107 34645 3135 34679
rect 3173 34645 3175 34679
rect 3175 34645 3207 34679
rect 3245 34645 3277 34679
rect 3277 34645 3279 34679
rect 3317 34645 3345 34679
rect 3345 34645 3351 34679
rect 3389 34645 3413 34679
rect 3413 34645 3423 34679
rect 3461 34645 3481 34679
rect 3481 34645 3495 34679
rect 3533 34645 3549 34679
rect 3549 34645 3567 34679
rect 3605 34645 3617 34679
rect 3617 34645 3639 34679
rect 3677 34645 3685 34679
rect 3685 34645 3711 34679
rect 3749 34645 3753 34679
rect 3753 34645 3783 34679
rect 3821 34645 3855 34679
rect 3893 34645 3923 34679
rect 3923 34645 3927 34679
rect 3965 34645 3991 34679
rect 3991 34645 3999 34679
rect 4037 34645 4059 34679
rect 4059 34645 4071 34679
rect 4109 34645 4127 34679
rect 4127 34645 4143 34679
rect 4181 34645 4195 34679
rect 4195 34645 4215 34679
rect 4253 34645 4263 34679
rect 4263 34645 4287 34679
rect 4325 34645 4331 34679
rect 4331 34645 4359 34679
rect 4397 34645 4399 34679
rect 4399 34645 4431 34679
rect 4469 34645 4501 34679
rect 4501 34645 4503 34679
rect 4541 34645 4569 34679
rect 4569 34645 4575 34679
rect 4613 34645 4637 34679
rect 4637 34645 4647 34679
rect 4685 34645 4705 34679
rect 4705 34645 4719 34679
rect 4757 34645 4773 34679
rect 4773 34645 4791 34679
rect 4829 34645 4841 34679
rect 4841 34645 4863 34679
rect 4901 34645 4909 34679
rect 4909 34645 4935 34679
rect 4973 34645 4977 34679
rect 4977 34645 5007 34679
rect 5045 34645 5079 34679
rect 5117 34645 5147 34679
rect 5147 34645 5151 34679
rect 5189 34645 5215 34679
rect 5215 34645 5223 34679
rect 5261 34645 5283 34679
rect 5283 34645 5295 34679
rect 5333 34645 5351 34679
rect 5351 34645 5367 34679
rect 5405 34645 5419 34679
rect 5419 34645 5439 34679
rect 5477 34645 5487 34679
rect 5487 34645 5511 34679
rect 5549 34645 5555 34679
rect 5555 34645 5583 34679
rect 5621 34645 5623 34679
rect 5623 34645 5655 34679
rect 5693 34645 5725 34679
rect 5725 34645 5727 34679
rect 5765 34645 5793 34679
rect 5793 34645 5799 34679
rect 5837 34645 5861 34679
rect 5861 34645 5871 34679
rect 5909 34645 5929 34679
rect 5929 34645 5943 34679
rect 5981 34645 5997 34679
rect 5997 34645 6015 34679
rect 6053 34645 6065 34679
rect 6065 34645 6087 34679
rect 6125 34645 6133 34679
rect 6133 34645 6159 34679
rect 6197 34645 6201 34679
rect 6201 34645 6231 34679
rect 6269 34645 6303 34679
rect 6341 34645 6371 34679
rect 6371 34645 6375 34679
rect 6413 34645 6439 34679
rect 6439 34645 6447 34679
rect 6485 34645 6507 34679
rect 6507 34645 6519 34679
rect 6557 34645 6575 34679
rect 6575 34645 6591 34679
rect 6629 34645 6643 34679
rect 6643 34645 6663 34679
rect 6701 34645 6711 34679
rect 6711 34645 6735 34679
rect 6773 34645 6779 34679
rect 6779 34645 6807 34679
rect 6845 34645 6847 34679
rect 6847 34645 6879 34679
rect 6917 34645 6949 34679
rect 6949 34645 6951 34679
rect 6989 34645 7017 34679
rect 7017 34645 7023 34679
rect 7061 34645 7085 34679
rect 7085 34645 7095 34679
rect 7133 34645 7153 34679
rect 7153 34645 7167 34679
rect 7205 34645 7221 34679
rect 7221 34645 7239 34679
rect 7277 34645 7289 34679
rect 7289 34645 7311 34679
rect 7349 34645 7357 34679
rect 7357 34645 7383 34679
rect 7421 34645 7425 34679
rect 7425 34645 7455 34679
rect 7493 34645 7527 34679
rect 7565 34645 7595 34679
rect 7595 34645 7599 34679
rect 7637 34645 7663 34679
rect 7663 34645 7671 34679
rect 7709 34645 7731 34679
rect 7731 34645 7743 34679
rect 7781 34645 7799 34679
rect 7799 34645 7815 34679
rect 7853 34645 7867 34679
rect 7867 34645 7887 34679
rect 7925 34645 7935 34679
rect 7935 34645 7959 34679
rect 7997 34645 8003 34679
rect 8003 34645 8031 34679
rect 8069 34645 8071 34679
rect 8071 34645 8103 34679
rect 8141 34645 8173 34679
rect 8173 34645 8175 34679
rect 8213 34645 8241 34679
rect 8241 34645 8247 34679
rect 8285 34645 8309 34679
rect 8309 34645 8319 34679
rect 8357 34645 8377 34679
rect 8377 34645 8391 34679
rect 8429 34645 8445 34679
rect 8445 34645 8463 34679
rect 8501 34645 8513 34679
rect 8513 34645 8535 34679
rect 8573 34645 8581 34679
rect 8581 34645 8607 34679
rect 8645 34645 8649 34679
rect 8649 34645 8679 34679
rect 8717 34645 8751 34679
rect 8789 34645 8819 34679
rect 8819 34645 8823 34679
rect 8861 34645 8887 34679
rect 8887 34645 8895 34679
rect 8933 34645 8955 34679
rect 8955 34645 8967 34679
rect 9005 34645 9023 34679
rect 9023 34645 9039 34679
rect 9077 34645 9091 34679
rect 9091 34645 9111 34679
rect 9149 34645 9159 34679
rect 9159 34645 9183 34679
rect 9221 34645 9227 34679
rect 9227 34645 9255 34679
rect 9293 34645 9295 34679
rect 9295 34645 9327 34679
rect 9365 34645 9397 34679
rect 9397 34645 9399 34679
rect 9437 34645 9465 34679
rect 9465 34645 9471 34679
rect 9509 34645 9533 34679
rect 9533 34645 9543 34679
rect 9581 34645 9601 34679
rect 9601 34645 9615 34679
rect 9653 34645 9669 34679
rect 9669 34645 9687 34679
rect 9725 34645 9737 34679
rect 9737 34645 9759 34679
rect 9797 34645 9805 34679
rect 9805 34645 9831 34679
rect 9869 34645 9873 34679
rect 9873 34645 9903 34679
rect 9941 34645 9975 34679
rect 10013 34645 10043 34679
rect 10043 34645 10047 34679
rect 10085 34645 10111 34679
rect 10111 34645 10119 34679
rect 10157 34645 10179 34679
rect 10179 34645 10191 34679
rect 10229 34645 10247 34679
rect 10247 34645 10263 34679
rect 10301 34645 10315 34679
rect 10315 34645 10335 34679
rect 10373 34645 10383 34679
rect 10383 34645 10407 34679
rect 10445 34645 10451 34679
rect 10451 34645 10479 34679
rect 10517 34645 10519 34679
rect 10519 34645 10551 34679
rect 10589 34645 10621 34679
rect 10621 34645 10623 34679
rect 10661 34645 10689 34679
rect 10689 34645 10695 34679
rect 10733 34645 10757 34679
rect 10757 34645 10767 34679
rect 10805 34645 10825 34679
rect 10825 34645 10839 34679
rect 10877 34645 10893 34679
rect 10893 34645 10911 34679
rect 10949 34645 10961 34679
rect 10961 34645 10983 34679
rect 11021 34645 11029 34679
rect 11029 34645 11055 34679
rect 11093 34645 11097 34679
rect 11097 34645 11127 34679
rect 11165 34645 11199 34679
rect 11237 34645 11267 34679
rect 11267 34645 11271 34679
rect 11309 34645 11335 34679
rect 11335 34645 11343 34679
rect 11381 34645 11403 34679
rect 11403 34645 11415 34679
rect 11453 34645 11471 34679
rect 11471 34645 11487 34679
rect 11525 34645 11539 34679
rect 11539 34645 11559 34679
rect 11597 34645 11607 34679
rect 11607 34645 11631 34679
rect 11669 34645 11675 34679
rect 11675 34645 11703 34679
rect 11741 34645 11743 34679
rect 11743 34645 11775 34679
rect 11813 34645 11845 34679
rect 11845 34645 11847 34679
rect 11885 34645 11913 34679
rect 11913 34645 11919 34679
rect 11957 34645 11981 34679
rect 11981 34645 11991 34679
rect 12029 34645 12049 34679
rect 12049 34645 12063 34679
rect 12101 34645 12117 34679
rect 12117 34645 12135 34679
rect 12173 34645 12185 34679
rect 12185 34645 12207 34679
rect 12245 34645 12253 34679
rect 12253 34645 12279 34679
rect 12317 34645 12321 34679
rect 12321 34645 12351 34679
rect 12389 34645 12423 34679
rect 12461 34645 12491 34679
rect 12491 34645 12495 34679
rect 12533 34645 12559 34679
rect 12559 34645 12567 34679
rect 12605 34645 12627 34679
rect 12627 34645 12639 34679
rect 12677 34645 12695 34679
rect 12695 34645 12711 34679
rect 12749 34645 12763 34679
rect 12763 34645 12783 34679
rect 12821 34645 12831 34679
rect 12831 34645 12855 34679
rect 12893 34645 12899 34679
rect 12899 34645 12927 34679
rect 12965 34645 12967 34679
rect 12967 34645 12999 34679
rect 13037 34645 13069 34679
rect 13069 34645 13071 34679
rect 13109 34645 13137 34679
rect 13137 34645 13143 34679
rect 13181 34645 13205 34679
rect 13205 34645 13215 34679
rect 13253 34645 13273 34679
rect 13273 34645 13287 34679
rect 13325 34645 13341 34679
rect 13341 34645 13359 34679
rect 13397 34645 13409 34679
rect 13409 34645 13431 34679
rect 13469 34645 13477 34679
rect 13477 34645 13503 34679
rect 13541 34645 13545 34679
rect 13545 34645 13575 34679
rect 13613 34645 13647 34679
rect 13685 34645 13715 34679
rect 13715 34645 13719 34679
rect 1161 34462 1195 34482
rect 1161 34448 1195 34462
rect 1161 34394 1195 34410
rect 1161 34376 1195 34394
rect 1161 34326 1195 34338
rect 1161 34304 1195 34326
rect 1161 34258 1195 34266
rect 1161 34232 1195 34258
rect 1161 34190 1195 34194
rect 1161 34160 1195 34190
rect 1161 34088 1195 34122
rect 1161 34020 1195 34050
rect 1161 34016 1195 34020
rect 1161 33952 1195 33978
rect 1161 33944 1195 33952
rect 1161 33884 1195 33906
rect 1161 33872 1195 33884
rect 1161 33816 1195 33834
rect 1161 33800 1195 33816
rect 1161 33748 1195 33762
rect 1161 33728 1195 33748
rect 1161 33680 1195 33690
rect 1161 33656 1195 33680
rect 1161 33612 1195 33618
rect 1161 33584 1195 33612
rect 1161 33544 1195 33546
rect 1161 33512 1195 33544
rect 1161 33442 1195 33474
rect 1161 33440 1195 33442
rect 1161 33374 1195 33402
rect 1161 33368 1195 33374
rect 1161 33306 1195 33330
rect 1161 33296 1195 33306
rect 1161 33238 1195 33258
rect 1161 33224 1195 33238
rect 1161 33170 1195 33186
rect 1161 33152 1195 33170
rect 1161 33102 1195 33114
rect 1161 33080 1195 33102
rect 1161 33034 1195 33042
rect 1161 33008 1195 33034
rect 1161 32966 1195 32970
rect 1161 32936 1195 32966
rect 1161 32864 1195 32898
rect 1161 32796 1195 32826
rect 1161 32792 1195 32796
rect 1161 32728 1195 32754
rect 1161 32720 1195 32728
rect 1161 32660 1195 32682
rect 1161 32648 1195 32660
rect 1161 32592 1195 32610
rect 1161 32576 1195 32592
rect 1161 32524 1195 32538
rect 1161 32504 1195 32524
rect 1161 32456 1195 32466
rect 1161 32432 1195 32456
rect 1161 32388 1195 32394
rect 1161 32360 1195 32388
rect 1161 32320 1195 32322
rect 1161 32288 1195 32320
rect 1161 32218 1195 32250
rect 1161 32216 1195 32218
rect 1161 32150 1195 32178
rect 1161 32144 1195 32150
rect 1161 32082 1195 32106
rect 1161 32072 1195 32082
rect 1161 32014 1195 32034
rect 1161 32000 1195 32014
rect 1161 31946 1195 31962
rect 1161 31928 1195 31946
rect 1161 31878 1195 31890
rect 1161 31856 1195 31878
rect 1161 31810 1195 31818
rect 1161 31784 1195 31810
rect 1161 31742 1195 31746
rect 1161 31712 1195 31742
rect 1161 31640 1195 31674
rect 1161 31572 1195 31602
rect 1161 31568 1195 31572
rect 1161 31504 1195 31530
rect 1161 31496 1195 31504
rect 1161 31436 1195 31458
rect 1161 31424 1195 31436
rect 1161 31368 1195 31386
rect 1161 31352 1195 31368
rect 1161 31300 1195 31314
rect 1161 31280 1195 31300
rect 1161 31232 1195 31242
rect 1161 31208 1195 31232
rect 1161 31164 1195 31170
rect 1161 31136 1195 31164
rect 1161 31096 1195 31098
rect 1161 31064 1195 31096
rect 1161 30994 1195 31026
rect 1161 30992 1195 30994
rect 1161 30926 1195 30954
rect 1161 30920 1195 30926
rect 1161 30858 1195 30882
rect 1161 30848 1195 30858
rect 1161 30790 1195 30810
rect 1161 30776 1195 30790
rect 1161 30722 1195 30738
rect 1161 30704 1195 30722
rect 1161 30654 1195 30666
rect 1161 30632 1195 30654
rect 1161 30586 1195 30594
rect 1161 30560 1195 30586
rect 1161 30518 1195 30522
rect 1161 30488 1195 30518
rect 1161 30416 1195 30450
rect 1161 30348 1195 30378
rect 1161 30344 1195 30348
rect 1161 30280 1195 30306
rect 1161 30272 1195 30280
rect 1161 30212 1195 30234
rect 1161 30200 1195 30212
rect 1161 30144 1195 30162
rect 1161 30128 1195 30144
rect 1161 30076 1195 30090
rect 1161 30056 1195 30076
rect 1161 30008 1195 30018
rect 1161 29984 1195 30008
rect 1161 29940 1195 29946
rect 1161 29912 1195 29940
rect 1161 29872 1195 29874
rect 1161 29840 1195 29872
rect 1161 29770 1195 29802
rect 1161 29768 1195 29770
rect 1161 29702 1195 29730
rect 1161 29696 1195 29702
rect 1161 29634 1195 29658
rect 1161 29624 1195 29634
rect 1161 29566 1195 29586
rect 1161 29552 1195 29566
rect 1161 29498 1195 29514
rect 1161 29480 1195 29498
rect 1161 29430 1195 29442
rect 1161 29408 1195 29430
rect 1161 29362 1195 29370
rect 1161 29336 1195 29362
rect 1161 29294 1195 29298
rect 1161 29264 1195 29294
rect 1161 29192 1195 29226
rect 1161 29124 1195 29154
rect 1161 29120 1195 29124
rect 1161 29056 1195 29082
rect 1161 29048 1195 29056
rect 1161 28988 1195 29010
rect 1161 28976 1195 28988
rect 1161 28920 1195 28938
rect 1161 28904 1195 28920
rect 13809 34457 13843 34474
rect 13809 34440 13843 34457
rect 13809 34389 13843 34402
rect 13809 34368 13843 34389
rect 13809 34321 13843 34330
rect 13809 34296 13843 34321
rect 13809 34253 13843 34258
rect 13809 34224 13843 34253
rect 13809 34185 13843 34186
rect 13809 34152 13843 34185
rect 13809 34083 13843 34114
rect 13809 34080 13843 34083
rect 13809 34015 13843 34042
rect 13809 34008 13843 34015
rect 13809 33947 13843 33970
rect 13809 33936 13843 33947
rect 13809 33879 13843 33898
rect 13809 33864 13843 33879
rect 13809 33811 13843 33826
rect 13809 33792 13843 33811
rect 13809 33743 13843 33754
rect 13809 33720 13843 33743
rect 13809 33675 13843 33682
rect 13809 33648 13843 33675
rect 13809 33607 13843 33610
rect 13809 33576 13843 33607
rect 13809 33505 13843 33538
rect 13809 33504 13843 33505
rect 13809 33437 13843 33466
rect 13809 33432 13843 33437
rect 13809 33369 13843 33394
rect 13809 33360 13843 33369
rect 13809 33301 13843 33322
rect 13809 33288 13843 33301
rect 13809 33233 13843 33250
rect 13809 33216 13843 33233
rect 13809 33165 13843 33178
rect 13809 33144 13843 33165
rect 13809 33097 13843 33106
rect 13809 33072 13843 33097
rect 13809 33029 13843 33034
rect 13809 33000 13843 33029
rect 13809 32961 13843 32962
rect 13809 32928 13843 32961
rect 13809 32859 13843 32890
rect 13809 32856 13843 32859
rect 13809 32791 13843 32818
rect 13809 32784 13843 32791
rect 13809 32723 13843 32746
rect 13809 32712 13843 32723
rect 13809 32655 13843 32674
rect 13809 32640 13843 32655
rect 13809 32587 13843 32602
rect 13809 32568 13843 32587
rect 13809 32519 13843 32530
rect 13809 32496 13843 32519
rect 13809 32451 13843 32458
rect 13809 32424 13843 32451
rect 13809 32383 13843 32386
rect 13809 32352 13843 32383
rect 13809 32281 13843 32314
rect 13809 32280 13843 32281
rect 13809 32213 13843 32242
rect 13809 32208 13843 32213
rect 13809 32145 13843 32170
rect 13809 32136 13843 32145
rect 13809 32077 13843 32098
rect 13809 32064 13843 32077
rect 13809 32009 13843 32026
rect 13809 31992 13843 32009
rect 13809 31941 13843 31954
rect 13809 31920 13843 31941
rect 13809 31873 13843 31882
rect 13809 31848 13843 31873
rect 13809 31805 13843 31810
rect 13809 31776 13843 31805
rect 13809 31737 13843 31738
rect 13809 31704 13843 31737
rect 13809 31635 13843 31666
rect 13809 31632 13843 31635
rect 13809 31567 13843 31594
rect 13809 31560 13843 31567
rect 13809 31499 13843 31522
rect 13809 31488 13843 31499
rect 13809 31431 13843 31450
rect 13809 31416 13843 31431
rect 13809 31363 13843 31378
rect 13809 31344 13843 31363
rect 13809 31295 13843 31306
rect 13809 31272 13843 31295
rect 13809 31227 13843 31234
rect 13809 31200 13843 31227
rect 13809 31159 13843 31162
rect 13809 31128 13843 31159
rect 13809 31057 13843 31090
rect 13809 31056 13843 31057
rect 13809 30989 13843 31018
rect 13809 30984 13843 30989
rect 13809 30921 13843 30946
rect 13809 30912 13843 30921
rect 13809 30853 13843 30874
rect 13809 30840 13843 30853
rect 13809 30785 13843 30802
rect 13809 30768 13843 30785
rect 13809 30717 13843 30730
rect 13809 30696 13843 30717
rect 13809 30649 13843 30658
rect 13809 30624 13843 30649
rect 13809 30581 13843 30586
rect 13809 30552 13843 30581
rect 13809 30513 13843 30514
rect 13809 30480 13843 30513
rect 13809 30411 13843 30442
rect 13809 30408 13843 30411
rect 13809 30343 13843 30370
rect 13809 30336 13843 30343
rect 13809 30275 13843 30298
rect 13809 30264 13843 30275
rect 13809 30207 13843 30226
rect 13809 30192 13843 30207
rect 13809 30139 13843 30154
rect 13809 30120 13843 30139
rect 13809 30071 13843 30082
rect 13809 30048 13843 30071
rect 13809 30003 13843 30010
rect 13809 29976 13843 30003
rect 13809 29935 13843 29938
rect 13809 29904 13843 29935
rect 13809 29833 13843 29866
rect 13809 29832 13843 29833
rect 13809 29765 13843 29794
rect 13809 29760 13843 29765
rect 13809 29697 13843 29722
rect 13809 29688 13843 29697
rect 13809 29629 13843 29650
rect 13809 29616 13843 29629
rect 13809 29561 13843 29578
rect 13809 29544 13843 29561
rect 13809 29493 13843 29506
rect 13809 29472 13843 29493
rect 13809 29425 13843 29434
rect 13809 29400 13843 29425
rect 13809 29357 13843 29362
rect 13809 29328 13843 29357
rect 13809 29289 13843 29290
rect 13809 29256 13843 29289
rect 13809 29187 13843 29218
rect 13809 29184 13843 29187
rect 13809 29119 13843 29146
rect 13809 29112 13843 29119
rect 13809 29051 13843 29074
rect 13809 29040 13843 29051
rect 13809 28983 13843 29002
rect 13809 28968 13843 28983
rect 1161 28852 1195 28866
rect 1161 28832 1195 28852
rect 1161 28784 1195 28794
rect 1161 28760 1195 28784
rect 1161 28716 1195 28722
rect 1161 28688 1195 28716
rect 1161 28648 1195 28650
rect 1161 28616 1195 28648
rect 1161 28546 1195 28578
rect 1161 28544 1195 28546
rect 1161 28478 1195 28506
rect 1161 28472 1195 28478
rect 1161 28410 1195 28434
rect 1161 28400 1195 28410
rect 1161 28342 1195 28362
rect 1161 28328 1195 28342
rect 1161 28274 1195 28290
rect 1161 28256 1195 28274
rect 1161 28206 1195 28218
rect 1161 28184 1195 28206
rect 1161 28138 1195 28146
rect 1161 28112 1195 28138
rect 1161 28070 1195 28074
rect 1161 28040 1195 28070
rect 1161 27968 1195 28002
rect 1161 27900 1195 27930
rect 1161 27896 1195 27900
rect 1161 27832 1195 27858
rect 1161 27824 1195 27832
rect 1161 27764 1195 27786
rect 1161 27752 1195 27764
rect 1161 27696 1195 27714
rect 1161 27680 1195 27696
rect 1161 27628 1195 27642
rect 1161 27608 1195 27628
rect 1161 27560 1195 27570
rect 1161 27536 1195 27560
rect 1161 27492 1195 27498
rect 1161 27464 1195 27492
rect 1161 27424 1195 27426
rect 1161 27392 1195 27424
rect 1161 27322 1195 27354
rect 1161 27320 1195 27322
rect 1161 27254 1195 27282
rect 1161 27248 1195 27254
rect 1161 27186 1195 27210
rect 1161 27176 1195 27186
rect 1161 27118 1195 27138
rect 1161 27104 1195 27118
rect 1161 27050 1195 27066
rect 1161 27032 1195 27050
rect 1982 28553 2119 28875
rect 2119 28553 12897 28875
rect 12897 28553 13032 28875
rect 1726 28422 1976 28489
rect 1726 27504 1976 28422
rect 13031 28422 13281 28482
rect 1726 27447 1976 27504
rect 13031 27504 13281 28422
rect 13031 27440 13281 27504
rect 1985 27084 2119 27334
rect 2119 27084 12897 27334
rect 12897 27084 13035 27334
rect 13809 28915 13843 28930
rect 13809 28896 13843 28915
rect 13809 28847 13843 28858
rect 13809 28824 13843 28847
rect 13809 28779 13843 28786
rect 13809 28752 13843 28779
rect 1161 26982 1195 26994
rect 1161 26960 1195 26982
rect 1161 26914 1195 26922
rect 1161 26888 1195 26914
rect 1161 26846 1195 26850
rect 1161 26816 1195 26846
rect 1161 26744 1195 26778
rect 1161 26676 1195 26706
rect 1161 26672 1195 26676
rect 1161 26608 1195 26634
rect 1161 26600 1195 26608
rect 1161 26540 1195 26562
rect 1161 26528 1195 26540
rect 1161 26472 1195 26490
rect 1161 26456 1195 26472
rect 1161 26404 1195 26418
rect 1161 26384 1195 26404
rect 1161 26336 1195 26346
rect 1161 26312 1195 26336
rect 1161 26268 1195 26274
rect 1161 26240 1195 26268
rect 1161 26200 1195 26202
rect 1161 26168 1195 26200
rect 1161 26098 1195 26130
rect 1161 26096 1195 26098
rect 1161 26030 1195 26058
rect 1161 26024 1195 26030
rect 1161 25962 1195 25986
rect 1161 25952 1195 25962
rect 1161 25894 1195 25914
rect 1161 25880 1195 25894
rect 1161 25826 1195 25842
rect 1161 25808 1195 25826
rect 1161 25758 1195 25770
rect 1161 25736 1195 25758
rect 1161 25690 1195 25698
rect 1161 25664 1195 25690
rect 1161 25622 1195 25626
rect 1161 25592 1195 25622
rect 1161 25520 1195 25554
rect 1161 25452 1195 25482
rect 1161 25448 1195 25452
rect 1161 25384 1195 25410
rect 1161 25376 1195 25384
rect 1161 25316 1195 25338
rect 1161 25304 1195 25316
rect 1161 25248 1195 25266
rect 1161 25232 1195 25248
rect 1161 25180 1195 25194
rect 1161 25160 1195 25180
rect 1161 25112 1195 25122
rect 1161 25088 1195 25112
rect 1161 25044 1195 25050
rect 1161 25016 1195 25044
rect 1161 24976 1195 24978
rect 1161 24944 1195 24976
rect 1161 24874 1195 24906
rect 1161 24872 1195 24874
rect 1161 24806 1195 24834
rect 1161 24800 1195 24806
rect 1161 24738 1195 24762
rect 1161 24728 1195 24738
rect 1161 24670 1195 24690
rect 1161 24656 1195 24670
rect 1161 24602 1195 24618
rect 1161 24584 1195 24602
rect 1161 24534 1195 24546
rect 1161 24512 1195 24534
rect 1161 24466 1195 24474
rect 1161 24440 1195 24466
rect 1161 24398 1195 24402
rect 1161 24368 1195 24398
rect 1161 24296 1195 24330
rect 1161 24228 1195 24258
rect 1161 24224 1195 24228
rect 1161 24160 1195 24186
rect 1161 24152 1195 24160
rect 1161 24092 1195 24114
rect 1161 24080 1195 24092
rect 1161 24024 1195 24042
rect 1161 24008 1195 24024
rect 1161 23956 1195 23970
rect 1161 23936 1195 23956
rect 1161 23888 1195 23898
rect 1161 23864 1195 23888
rect 1161 23820 1195 23826
rect 1161 23792 1195 23820
rect 1161 23752 1195 23754
rect 1161 23720 1195 23752
rect 1161 23650 1195 23682
rect 1161 23648 1195 23650
rect 1161 23582 1195 23610
rect 1161 23576 1195 23582
rect 1161 23514 1195 23538
rect 1161 23504 1195 23514
rect 1161 23446 1195 23466
rect 1161 23432 1195 23446
rect 1161 23378 1195 23394
rect 1161 23360 1195 23378
rect 1161 23310 1195 23322
rect 1161 23288 1195 23310
rect 1161 23242 1195 23250
rect 1161 23216 1195 23242
rect 1161 23174 1195 23178
rect 1161 23144 1195 23174
rect 1161 23072 1195 23106
rect 1161 23004 1195 23034
rect 1161 23000 1195 23004
rect 1161 22936 1195 22962
rect 1161 22928 1195 22936
rect 1161 22868 1195 22890
rect 1161 22856 1195 22868
rect 1161 22800 1195 22818
rect 1161 22784 1195 22800
rect 1161 22732 1195 22746
rect 1161 22712 1195 22732
rect 1161 22664 1195 22674
rect 1161 22640 1195 22664
rect 1161 22596 1195 22602
rect 1161 22568 1195 22596
rect 1161 22528 1195 22530
rect 1161 22496 1195 22528
rect 1161 22426 1195 22458
rect 1161 22424 1195 22426
rect 1161 22358 1195 22386
rect 1161 22352 1195 22358
rect 1161 22290 1195 22314
rect 1161 22280 1195 22290
rect 1161 22222 1195 22242
rect 1161 22208 1195 22222
rect 1161 22154 1195 22170
rect 1161 22136 1195 22154
rect 1161 22086 1195 22098
rect 1161 22064 1195 22086
rect 1161 22018 1195 22026
rect 1161 21992 1195 22018
rect 1161 21950 1195 21954
rect 1161 21920 1195 21950
rect 1161 21848 1195 21882
rect 1161 21780 1195 21810
rect 1161 21776 1195 21780
rect 1161 21712 1195 21738
rect 1161 21704 1195 21712
rect 1161 21644 1195 21666
rect 1161 21632 1195 21644
rect 1161 21576 1195 21594
rect 1161 21560 1195 21576
rect 1161 21508 1195 21522
rect 1161 21488 1195 21508
rect 1161 21440 1195 21450
rect 1161 21416 1195 21440
rect 1161 21372 1195 21378
rect 1161 21344 1195 21372
rect 1161 21304 1195 21306
rect 1161 21272 1195 21304
rect 1161 21202 1195 21234
rect 1161 21200 1195 21202
rect 1161 21134 1195 21162
rect 1161 21128 1195 21134
rect 1161 21066 1195 21090
rect 1161 21056 1195 21066
rect 1161 20998 1195 21018
rect 1161 20984 1195 20998
rect 1161 20930 1195 20946
rect 1161 20912 1195 20930
rect 1161 20862 1195 20874
rect 1161 20840 1195 20862
rect 1161 20794 1195 20802
rect 1161 20768 1195 20794
rect 1161 20726 1195 20730
rect 1161 20696 1195 20726
rect 1161 20624 1195 20658
rect 1161 20556 1195 20586
rect 1161 20552 1195 20556
rect 1161 20488 1195 20514
rect 1161 20480 1195 20488
rect 1161 20420 1195 20442
rect 1161 20408 1195 20420
rect 1161 20352 1195 20370
rect 1161 20336 1195 20352
rect 1161 20284 1195 20298
rect 1161 20264 1195 20284
rect 1161 20216 1195 20226
rect 1161 20192 1195 20216
rect 1161 20148 1195 20154
rect 1161 20120 1195 20148
rect 1161 20080 1195 20082
rect 1161 20048 1195 20080
rect 1161 19978 1195 20010
rect 1161 19976 1195 19978
rect 1161 19910 1195 19938
rect 1161 19904 1195 19910
rect 1161 19842 1195 19866
rect 1161 19832 1195 19842
rect 1161 19774 1195 19794
rect 1161 19760 1195 19774
rect 1161 19706 1195 19722
rect 1161 19688 1195 19706
rect 1161 19638 1195 19650
rect 1161 19616 1195 19638
rect 1161 19570 1195 19578
rect 1161 19544 1195 19570
rect 1161 19502 1195 19506
rect 1161 19472 1195 19502
rect 1161 19400 1195 19434
rect 1161 19332 1195 19362
rect 1161 19328 1195 19332
rect 1161 19264 1195 19290
rect 1161 19256 1195 19264
rect 1161 19196 1195 19218
rect 1161 19184 1195 19196
rect 1161 19128 1195 19146
rect 1161 19112 1195 19128
rect 1161 19060 1195 19074
rect 1161 19040 1195 19060
rect 1161 18992 1195 19002
rect 1161 18968 1195 18992
rect 1161 18924 1195 18930
rect 1161 18896 1195 18924
rect 1161 18856 1195 18858
rect 1161 18824 1195 18856
rect 1161 18754 1195 18786
rect 1161 18752 1195 18754
rect 1161 18686 1195 18714
rect 1161 18680 1195 18686
rect 1161 18618 1195 18642
rect 1161 18608 1195 18618
rect 1161 18550 1195 18570
rect 1161 18536 1195 18550
rect 1161 18482 1195 18498
rect 1161 18464 1195 18482
rect 1161 18414 1195 18426
rect 1161 18392 1195 18414
rect 1161 18346 1195 18354
rect 1161 18320 1195 18346
rect 1161 18278 1195 18282
rect 1161 18248 1195 18278
rect 1161 18176 1195 18210
rect 1161 18108 1195 18138
rect 1161 18104 1195 18108
rect 1161 18040 1195 18066
rect 1161 18032 1195 18040
rect 1161 17972 1195 17994
rect 1161 17960 1195 17972
rect 1161 17904 1195 17922
rect 1161 17888 1195 17904
rect 1161 17836 1195 17850
rect 1161 17816 1195 17836
rect 1161 17768 1195 17778
rect 1161 17744 1195 17768
rect 1161 17700 1195 17706
rect 1161 17672 1195 17700
rect 1161 17632 1195 17634
rect 1161 17600 1195 17632
rect 1161 17530 1195 17562
rect 1161 17528 1195 17530
rect 1161 17462 1195 17490
rect 1161 17456 1195 17462
rect 1161 17394 1195 17418
rect 1161 17384 1195 17394
rect 1161 17326 1195 17346
rect 1161 17312 1195 17326
rect 1161 17258 1195 17274
rect 1161 17240 1195 17258
rect 1161 17190 1195 17202
rect 1161 17168 1195 17190
rect 1161 17122 1195 17130
rect 1161 17096 1195 17122
rect 1161 17054 1195 17058
rect 1161 17024 1195 17054
rect 1161 16952 1195 16986
rect 1161 16884 1195 16914
rect 1161 16880 1195 16884
rect 1161 16816 1195 16842
rect 1161 16808 1195 16816
rect 1161 16748 1195 16770
rect 1161 16736 1195 16748
rect 1161 16680 1195 16698
rect 1161 16664 1195 16680
rect 1161 16612 1195 16626
rect 1161 16592 1195 16612
rect 1161 16544 1195 16554
rect 1161 16520 1195 16544
rect 1161 16476 1195 16482
rect 1161 16448 1195 16476
rect 1161 16408 1195 16410
rect 1161 16376 1195 16408
rect 1161 16306 1195 16338
rect 1161 16304 1195 16306
rect 1161 16238 1195 16266
rect 1161 16232 1195 16238
rect 1161 16170 1195 16194
rect 1161 16160 1195 16170
rect 1161 16102 1195 16122
rect 1161 16088 1195 16102
rect 1161 16034 1195 16050
rect 1161 16016 1195 16034
rect 1161 15966 1195 15978
rect 1161 15944 1195 15966
rect 1161 15898 1195 15906
rect 1161 15872 1195 15898
rect 1161 15830 1195 15834
rect 1161 15800 1195 15830
rect 1161 15728 1195 15762
rect 1161 15660 1195 15690
rect 1161 15656 1195 15660
rect 1161 15592 1195 15618
rect 1161 15584 1195 15592
rect 1161 15524 1195 15546
rect 1161 15512 1195 15524
rect 1161 15456 1195 15474
rect 1161 15440 1195 15456
rect 1161 15388 1195 15402
rect 1161 15368 1195 15388
rect 13809 23373 13843 23397
rect 13809 23363 13843 23373
rect 13809 23305 13843 23325
rect 13809 23291 13843 23305
rect 13809 23237 13843 23253
rect 13809 23219 13843 23237
rect 13809 23169 13843 23181
rect 13809 23147 13843 23169
rect 13809 23101 13843 23109
rect 13809 23075 13843 23101
rect 13809 23033 13843 23037
rect 13809 23003 13843 23033
rect 13809 22931 13843 22965
rect 13809 22863 13843 22893
rect 13809 22859 13843 22863
rect 13809 22795 13843 22821
rect 13809 22787 13843 22795
rect 13809 22727 13843 22749
rect 13809 22715 13843 22727
rect 13809 22659 13843 22677
rect 13809 22643 13843 22659
rect 13809 22591 13843 22605
rect 13809 22571 13843 22591
rect 13809 22523 13843 22533
rect 13809 22499 13843 22523
rect 13809 22455 13843 22461
rect 13809 22427 13843 22455
rect 13809 22387 13843 22389
rect 13809 22355 13843 22387
rect 13809 22285 13843 22317
rect 13809 22283 13843 22285
rect 13809 22217 13843 22245
rect 13809 22211 13843 22217
rect 13809 22149 13843 22173
rect 13809 22139 13843 22149
rect 13809 22081 13843 22101
rect 13809 22067 13843 22081
rect 13809 22013 13843 22029
rect 13809 21995 13843 22013
rect 13809 21945 13843 21957
rect 13809 21923 13843 21945
rect 13809 21877 13843 21885
rect 13809 21851 13843 21877
rect 13809 21809 13843 21813
rect 13809 21779 13843 21809
rect 13809 21707 13843 21741
rect 13809 21639 13843 21669
rect 13809 21635 13843 21639
rect 13809 21571 13843 21597
rect 13809 21563 13843 21571
rect 13809 21503 13843 21525
rect 13809 21491 13843 21503
rect 13809 21435 13843 21453
rect 13809 21419 13843 21435
rect 13809 21367 13843 21381
rect 13809 21347 13843 21367
rect 13809 21299 13843 21309
rect 13809 21275 13843 21299
rect 13809 21231 13843 21237
rect 13809 21203 13843 21231
rect 13809 21163 13843 21165
rect 13809 21131 13843 21163
rect 13809 21061 13843 21093
rect 13809 21059 13843 21061
rect 13809 20993 13843 21021
rect 13809 20987 13843 20993
rect 13809 20925 13843 20949
rect 13809 20915 13843 20925
rect 13809 20857 13843 20877
rect 13809 20843 13843 20857
rect 13809 20789 13843 20805
rect 13809 20771 13843 20789
rect 13809 20721 13843 20733
rect 13809 20699 13843 20721
rect 13809 20653 13843 20661
rect 13809 20627 13843 20653
rect 13809 20585 13843 20589
rect 13809 20555 13843 20585
rect 13809 20483 13843 20517
rect 13809 20415 13843 20445
rect 13809 20411 13843 20415
rect 13809 20347 13843 20373
rect 13809 20339 13843 20347
rect 13809 20279 13843 20301
rect 13809 20267 13843 20279
rect 13809 20211 13843 20229
rect 13809 20195 13843 20211
rect 13809 20143 13843 20157
rect 13809 20123 13843 20143
rect 13809 20075 13843 20085
rect 13809 20051 13843 20075
rect 13809 20007 13843 20013
rect 13809 19979 13843 20007
rect 13809 19939 13843 19941
rect 13809 19907 13843 19939
rect 13809 19837 13843 19869
rect 13809 19835 13843 19837
rect 13809 19769 13843 19797
rect 13809 19763 13843 19769
rect 13809 19701 13843 19725
rect 13809 19691 13843 19701
rect 13809 19633 13843 19653
rect 13809 19619 13843 19633
rect 13809 19565 13843 19581
rect 13809 19547 13843 19565
rect 13809 19497 13843 19509
rect 13809 19475 13843 19497
rect 13809 19429 13843 19437
rect 13809 19403 13843 19429
rect 13809 19361 13843 19365
rect 13809 19331 13843 19361
rect 13809 19259 13843 19293
rect 13809 19191 13843 19221
rect 13809 19187 13843 19191
rect 13809 19123 13843 19149
rect 13809 19115 13843 19123
rect 13809 19055 13843 19077
rect 13809 19043 13843 19055
rect 13809 18987 13843 19005
rect 13809 18971 13843 18987
rect 13809 18919 13843 18933
rect 13809 18899 13843 18919
rect 13809 18851 13843 18861
rect 13809 18827 13843 18851
rect 13809 18783 13843 18789
rect 13809 18755 13843 18783
rect 13809 18715 13843 18717
rect 13809 18683 13843 18715
rect 13809 18613 13843 18645
rect 13809 18611 13843 18613
rect 13809 18545 13843 18573
rect 13809 18539 13843 18545
rect 13809 18477 13843 18501
rect 13809 18467 13843 18477
rect 13809 18409 13843 18429
rect 13809 18395 13843 18409
rect 13809 18341 13843 18357
rect 13809 18323 13843 18341
rect 13809 18273 13843 18285
rect 13809 18251 13843 18273
rect 13809 18205 13843 18213
rect 13809 18179 13843 18205
rect 13809 18137 13843 18141
rect 13809 18107 13843 18137
rect 13809 18035 13843 18069
rect 13809 17967 13843 17997
rect 13809 17963 13843 17967
rect 13809 17899 13843 17925
rect 13809 17891 13843 17899
rect 13809 17831 13843 17853
rect 13809 17819 13843 17831
rect 13809 17763 13843 17781
rect 13809 17747 13843 17763
rect 13809 17695 13843 17709
rect 13809 17675 13843 17695
rect 13809 17627 13843 17637
rect 13809 17603 13843 17627
rect 13809 17559 13843 17565
rect 13809 17531 13843 17559
rect 13809 17491 13843 17493
rect 13809 17459 13843 17491
rect 13809 17389 13843 17421
rect 13809 17387 13843 17389
rect 13809 17321 13843 17349
rect 13809 17315 13843 17321
rect 13809 17253 13843 17277
rect 13809 17243 13843 17253
rect 13809 17185 13843 17205
rect 13809 17171 13843 17185
rect 13809 17117 13843 17133
rect 13809 17099 13843 17117
rect 13809 17049 13843 17061
rect 13809 17027 13843 17049
rect 13809 16981 13843 16989
rect 13809 16955 13843 16981
rect 13809 16913 13843 16917
rect 13809 16883 13843 16913
rect 13809 16811 13843 16845
rect 13809 16743 13843 16773
rect 13809 16739 13843 16743
rect 13809 16675 13843 16701
rect 13809 16667 13843 16675
rect 13809 16607 13843 16629
rect 13809 16595 13843 16607
rect 13809 16539 13843 16557
rect 13809 16523 13843 16539
rect 13809 16471 13843 16485
rect 13809 16451 13843 16471
rect 13809 16403 13843 16413
rect 13809 16379 13843 16403
rect 13809 16335 13843 16341
rect 13809 16307 13843 16335
rect 13809 16267 13843 16269
rect 13809 16235 13843 16267
rect 13809 16165 13843 16197
rect 13809 16163 13843 16165
rect 13809 16097 13843 16125
rect 13809 16091 13843 16097
rect 13809 16029 13843 16053
rect 13809 16019 13843 16029
rect 13809 15961 13843 15981
rect 13809 15947 13843 15961
rect 13809 15893 13843 15909
rect 13809 15875 13843 15893
rect 13809 15825 13843 15837
rect 13809 15803 13843 15825
rect 13809 15757 13843 15765
rect 13809 15731 13843 15757
rect 13809 15689 13843 15693
rect 13809 15659 13843 15689
rect 13809 15587 13843 15621
rect 13809 15519 13843 15549
rect 13809 15515 13843 15519
rect 13809 15451 13843 15477
rect 13809 15443 13843 15451
rect 13809 15383 13843 15405
rect 13809 15371 13843 15383
rect 1298 15244 1302 15278
rect 1302 15244 1332 15278
rect 1370 15244 1404 15278
rect 1442 15244 1472 15278
rect 1472 15244 1476 15278
rect 1514 15244 1540 15278
rect 1540 15244 1548 15278
rect 1586 15244 1608 15278
rect 1608 15244 1620 15278
rect 1658 15244 1676 15278
rect 1676 15244 1692 15278
rect 1730 15244 1744 15278
rect 1744 15244 1764 15278
rect 1802 15244 1812 15278
rect 1812 15244 1836 15278
rect 1874 15244 1880 15278
rect 1880 15244 1908 15278
rect 1946 15244 1948 15278
rect 1948 15244 1980 15278
rect 2018 15244 2050 15278
rect 2050 15244 2052 15278
rect 2090 15244 2118 15278
rect 2118 15244 2124 15278
rect 2162 15244 2186 15278
rect 2186 15244 2196 15278
rect 2234 15244 2254 15278
rect 2254 15244 2268 15278
rect 2306 15244 2322 15278
rect 2322 15244 2340 15278
rect 2378 15244 2390 15278
rect 2390 15244 2412 15278
rect 2450 15244 2458 15278
rect 2458 15244 2484 15278
rect 2522 15244 2526 15278
rect 2526 15244 2556 15278
rect 2594 15244 2628 15278
rect 2666 15244 2696 15278
rect 2696 15244 2700 15278
rect 2738 15244 2764 15278
rect 2764 15244 2772 15278
rect 2810 15244 2832 15278
rect 2832 15244 2844 15278
rect 2882 15244 2900 15278
rect 2900 15244 2916 15278
rect 2954 15244 2968 15278
rect 2968 15244 2988 15278
rect 3026 15244 3036 15278
rect 3036 15244 3060 15278
rect 3098 15244 3104 15278
rect 3104 15244 3132 15278
rect 3170 15244 3172 15278
rect 3172 15244 3204 15278
rect 3242 15244 3274 15278
rect 3274 15244 3276 15278
rect 3314 15244 3342 15278
rect 3342 15244 3348 15278
rect 3386 15244 3410 15278
rect 3410 15244 3420 15278
rect 3458 15244 3478 15278
rect 3478 15244 3492 15278
rect 3530 15244 3546 15278
rect 3546 15244 3564 15278
rect 3602 15244 3614 15278
rect 3614 15244 3636 15278
rect 3674 15244 3682 15278
rect 3682 15244 3708 15278
rect 3746 15244 3750 15278
rect 3750 15244 3780 15278
rect 3818 15244 3852 15278
rect 3890 15244 3920 15278
rect 3920 15244 3924 15278
rect 3962 15244 3988 15278
rect 3988 15244 3996 15278
rect 4034 15244 4056 15278
rect 4056 15244 4068 15278
rect 4106 15244 4124 15278
rect 4124 15244 4140 15278
rect 4178 15244 4192 15278
rect 4192 15244 4212 15278
rect 4250 15244 4260 15278
rect 4260 15244 4284 15278
rect 4322 15244 4328 15278
rect 4328 15244 4356 15278
rect 4394 15244 4396 15278
rect 4396 15244 4428 15278
rect 4466 15244 4498 15278
rect 4498 15244 4500 15278
rect 4538 15244 4566 15278
rect 4566 15244 4572 15278
rect 4610 15244 4634 15278
rect 4634 15244 4644 15278
rect 4682 15244 4702 15278
rect 4702 15244 4716 15278
rect 4754 15244 4770 15278
rect 4770 15244 4788 15278
rect 4826 15244 4838 15278
rect 4838 15244 4860 15278
rect 4898 15244 4906 15278
rect 4906 15244 4932 15278
rect 4970 15244 4974 15278
rect 4974 15244 5004 15278
rect 5042 15244 5076 15278
rect 5114 15244 5144 15278
rect 5144 15244 5148 15278
rect 5186 15244 5212 15278
rect 5212 15244 5220 15278
rect 5258 15244 5280 15278
rect 5280 15244 5292 15278
rect 5330 15244 5348 15278
rect 5348 15244 5364 15278
rect 5402 15244 5416 15278
rect 5416 15244 5436 15278
rect 5474 15244 5484 15278
rect 5484 15244 5508 15278
rect 5546 15244 5552 15278
rect 5552 15244 5580 15278
rect 5618 15244 5620 15278
rect 5620 15244 5652 15278
rect 5690 15244 5722 15278
rect 5722 15244 5724 15278
rect 5762 15244 5790 15278
rect 5790 15244 5796 15278
rect 5834 15244 5858 15278
rect 5858 15244 5868 15278
rect 5906 15244 5926 15278
rect 5926 15244 5940 15278
rect 5978 15244 5994 15278
rect 5994 15244 6012 15278
rect 6050 15244 6062 15278
rect 6062 15244 6084 15278
rect 6122 15244 6130 15278
rect 6130 15244 6156 15278
rect 6194 15244 6198 15278
rect 6198 15244 6228 15278
rect 6266 15244 6300 15278
rect 6338 15244 6368 15278
rect 6368 15244 6372 15278
rect 6410 15244 6436 15278
rect 6436 15244 6444 15278
rect 6482 15244 6504 15278
rect 6504 15244 6516 15278
rect 6554 15244 6572 15278
rect 6572 15244 6588 15278
rect 6626 15244 6640 15278
rect 6640 15244 6660 15278
rect 6698 15244 6708 15278
rect 6708 15244 6732 15278
rect 6770 15244 6776 15278
rect 6776 15244 6804 15278
rect 6842 15244 6844 15278
rect 6844 15244 6876 15278
rect 6914 15244 6946 15278
rect 6946 15244 6948 15278
rect 6986 15244 7014 15278
rect 7014 15244 7020 15278
rect 7058 15244 7082 15278
rect 7082 15244 7092 15278
rect 7130 15244 7150 15278
rect 7150 15244 7164 15278
rect 7202 15244 7218 15278
rect 7218 15244 7236 15278
rect 7274 15244 7286 15278
rect 7286 15244 7308 15278
rect 7346 15244 7354 15278
rect 7354 15244 7380 15278
rect 7418 15244 7422 15278
rect 7422 15244 7452 15278
rect 7490 15244 7524 15278
rect 7562 15244 7592 15278
rect 7592 15244 7596 15278
rect 7634 15244 7660 15278
rect 7660 15244 7668 15278
rect 7706 15244 7728 15278
rect 7728 15244 7740 15278
rect 7778 15244 7796 15278
rect 7796 15244 7812 15278
rect 7850 15244 7864 15278
rect 7864 15244 7884 15278
rect 7922 15244 7932 15278
rect 7932 15244 7956 15278
rect 7994 15244 8000 15278
rect 8000 15244 8028 15278
rect 8066 15244 8068 15278
rect 8068 15244 8100 15278
rect 8138 15244 8170 15278
rect 8170 15244 8172 15278
rect 8210 15244 8238 15278
rect 8238 15244 8244 15278
rect 8282 15244 8306 15278
rect 8306 15244 8316 15278
rect 8354 15244 8374 15278
rect 8374 15244 8388 15278
rect 8426 15244 8442 15278
rect 8442 15244 8460 15278
rect 8498 15244 8510 15278
rect 8510 15244 8532 15278
rect 8570 15244 8578 15278
rect 8578 15244 8604 15278
rect 8642 15244 8646 15278
rect 8646 15244 8676 15278
rect 8714 15244 8748 15278
rect 8786 15244 8816 15278
rect 8816 15244 8820 15278
rect 8858 15244 8884 15278
rect 8884 15244 8892 15278
rect 8930 15244 8952 15278
rect 8952 15244 8964 15278
rect 9002 15244 9020 15278
rect 9020 15244 9036 15278
rect 9074 15244 9088 15278
rect 9088 15244 9108 15278
rect 9146 15244 9156 15278
rect 9156 15244 9180 15278
rect 9218 15244 9224 15278
rect 9224 15244 9252 15278
rect 9290 15244 9292 15278
rect 9292 15244 9324 15278
rect 9362 15244 9394 15278
rect 9394 15244 9396 15278
rect 9434 15244 9462 15278
rect 9462 15244 9468 15278
rect 9506 15244 9530 15278
rect 9530 15244 9540 15278
rect 9578 15244 9598 15278
rect 9598 15244 9612 15278
rect 9650 15244 9666 15278
rect 9666 15244 9684 15278
rect 9722 15244 9734 15278
rect 9734 15244 9756 15278
rect 9794 15244 9802 15278
rect 9802 15244 9828 15278
rect 9866 15244 9870 15278
rect 9870 15244 9900 15278
rect 9938 15244 9972 15278
rect 10010 15244 10040 15278
rect 10040 15244 10044 15278
rect 10082 15244 10108 15278
rect 10108 15244 10116 15278
rect 10154 15244 10176 15278
rect 10176 15244 10188 15278
rect 10226 15244 10244 15278
rect 10244 15244 10260 15278
rect 10298 15244 10312 15278
rect 10312 15244 10332 15278
rect 10370 15244 10380 15278
rect 10380 15244 10404 15278
rect 10442 15244 10448 15278
rect 10448 15244 10476 15278
rect 10514 15244 10516 15278
rect 10516 15244 10548 15278
rect 10586 15244 10618 15278
rect 10618 15244 10620 15278
rect 10658 15244 10686 15278
rect 10686 15244 10692 15278
rect 10730 15244 10754 15278
rect 10754 15244 10764 15278
rect 10802 15244 10822 15278
rect 10822 15244 10836 15278
rect 10874 15244 10890 15278
rect 10890 15244 10908 15278
rect 10946 15244 10958 15278
rect 10958 15244 10980 15278
rect 11018 15244 11026 15278
rect 11026 15244 11052 15278
rect 11090 15244 11094 15278
rect 11094 15244 11124 15278
rect 11162 15244 11196 15278
rect 11234 15244 11264 15278
rect 11264 15244 11268 15278
rect 11306 15244 11332 15278
rect 11332 15244 11340 15278
rect 11378 15244 11400 15278
rect 11400 15244 11412 15278
rect 11450 15244 11468 15278
rect 11468 15244 11484 15278
rect 11522 15244 11536 15278
rect 11536 15244 11556 15278
rect 11594 15244 11604 15278
rect 11604 15244 11628 15278
rect 11666 15244 11672 15278
rect 11672 15244 11700 15278
rect 11738 15244 11740 15278
rect 11740 15244 11772 15278
rect 11810 15244 11842 15278
rect 11842 15244 11844 15278
rect 11882 15244 11910 15278
rect 11910 15244 11916 15278
rect 11954 15244 11978 15278
rect 11978 15244 11988 15278
rect 12026 15244 12046 15278
rect 12046 15244 12060 15278
rect 12098 15244 12114 15278
rect 12114 15244 12132 15278
rect 12170 15244 12182 15278
rect 12182 15244 12204 15278
rect 12242 15244 12250 15278
rect 12250 15244 12276 15278
rect 12314 15244 12318 15278
rect 12318 15244 12348 15278
rect 12386 15244 12420 15278
rect 12458 15244 12488 15278
rect 12488 15244 12492 15278
rect 12530 15244 12556 15278
rect 12556 15244 12564 15278
rect 12602 15244 12624 15278
rect 12624 15244 12636 15278
rect 12674 15244 12692 15278
rect 12692 15244 12708 15278
rect 12746 15244 12760 15278
rect 12760 15244 12780 15278
rect 12818 15244 12828 15278
rect 12828 15244 12852 15278
rect 12890 15244 12896 15278
rect 12896 15244 12924 15278
rect 12962 15244 12964 15278
rect 12964 15244 12996 15278
rect 13034 15244 13066 15278
rect 13066 15244 13068 15278
rect 13106 15244 13134 15278
rect 13134 15244 13140 15278
rect 13178 15244 13202 15278
rect 13202 15244 13212 15278
rect 13250 15244 13270 15278
rect 13270 15244 13284 15278
rect 13322 15244 13338 15278
rect 13338 15244 13356 15278
rect 13394 15244 13406 15278
rect 13406 15244 13428 15278
rect 13466 15244 13474 15278
rect 13474 15244 13500 15278
rect 13538 15244 13542 15278
rect 13542 15244 13572 15278
rect 13610 15244 13644 15278
rect 13682 15244 13712 15278
rect 13712 15244 13716 15278
rect 14122 34707 14156 34741
rect 14122 34635 14156 34669
rect 14122 34563 14156 34597
rect 14122 34491 14156 34525
rect 14122 34419 14156 34453
rect 14122 34347 14156 34381
rect 14122 34275 14156 34309
rect 14122 34203 14156 34237
rect 14122 34131 14156 34165
rect 14122 34059 14156 34093
rect 14122 33987 14156 34021
rect 14122 33915 14156 33949
rect 14122 33843 14156 33877
rect 14122 33771 14156 33805
rect 14122 33699 14156 33733
rect 14122 33627 14156 33661
rect 14122 33555 14156 33589
rect 14122 33483 14156 33517
rect 14122 33411 14156 33445
rect 14122 33339 14156 33373
rect 14122 33267 14156 33301
rect 14122 33195 14156 33229
rect 14122 33123 14156 33157
rect 14122 33051 14156 33085
rect 14122 32979 14156 33013
rect 14122 32907 14156 32941
rect 14122 32835 14156 32869
rect 14122 32763 14156 32797
rect 14122 32691 14156 32725
rect 14122 32619 14156 32653
rect 14122 32547 14156 32581
rect 14122 32475 14156 32509
rect 14122 32403 14156 32437
rect 14122 32331 14156 32365
rect 14122 32259 14156 32293
rect 14122 32187 14156 32221
rect 14122 32115 14156 32149
rect 14122 32043 14156 32077
rect 14122 31971 14156 32005
rect 14122 31899 14156 31933
rect 14122 31827 14156 31861
rect 14122 31755 14156 31789
rect 14122 31683 14156 31717
rect 14122 31611 14156 31645
rect 14122 31539 14156 31573
rect 14122 31467 14156 31501
rect 14122 31395 14156 31429
rect 14122 31323 14156 31357
rect 14122 31251 14156 31285
rect 14122 31179 14156 31213
rect 14122 31107 14156 31141
rect 14122 31035 14156 31069
rect 14122 30963 14156 30997
rect 14122 30891 14156 30925
rect 14122 30819 14156 30853
rect 14122 30747 14156 30781
rect 14122 30675 14156 30709
rect 14122 30603 14156 30637
rect 14122 30531 14156 30565
rect 14122 30459 14156 30493
rect 14122 30387 14156 30421
rect 14122 30315 14156 30349
rect 14122 30243 14156 30277
rect 14122 30171 14156 30205
rect 14122 30099 14156 30133
rect 14122 30027 14156 30061
rect 14122 29955 14156 29989
rect 14122 29883 14156 29917
rect 14122 29811 14156 29845
rect 14122 29739 14156 29773
rect 14122 29667 14156 29701
rect 14122 29595 14156 29629
rect 14122 29523 14156 29557
rect 14122 29451 14156 29485
rect 14122 29379 14156 29413
rect 14122 29307 14156 29341
rect 14122 29235 14156 29269
rect 14122 29163 14156 29197
rect 14122 29091 14156 29125
rect 14122 29019 14156 29053
rect 14122 28947 14156 28981
rect 14122 28875 14156 28909
rect 14122 28803 14156 28837
rect 14122 28731 14156 28765
rect 14122 28659 14156 28693
rect 14122 28587 14156 28621
rect 14122 28515 14156 28549
rect 14122 28443 14156 28477
rect 14122 28371 14156 28405
rect 14122 28299 14156 28333
rect 14122 28227 14156 28261
rect 14122 28155 14156 28189
rect 14122 28083 14156 28117
rect 14122 28011 14156 28045
rect 14122 27939 14156 27973
rect 14122 27867 14156 27901
rect 14122 27795 14156 27829
rect 14122 27723 14156 27757
rect 14122 27651 14156 27685
rect 14122 27579 14156 27613
rect 14122 27507 14156 27541
rect 14122 27435 14156 27469
rect 14122 27363 14156 27397
rect 14122 27291 14156 27325
rect 14122 27219 14156 27253
rect 14122 27147 14156 27181
rect 14122 27075 14156 27109
rect 14122 27003 14156 27037
rect 14122 26931 14156 26965
rect 14122 26859 14156 26893
rect 14122 26787 14156 26821
rect 14122 26715 14156 26749
rect 14122 26643 14156 26677
rect 14122 26571 14156 26605
rect 14122 26499 14156 26533
rect 14122 26427 14156 26461
rect 14122 26355 14156 26389
rect 14122 26283 14156 26317
rect 14122 26211 14156 26245
rect 14122 26139 14156 26173
rect 14122 26067 14156 26101
rect 14122 25995 14156 26029
rect 14122 25923 14156 25957
rect 14122 25851 14156 25885
rect 14122 25779 14156 25813
rect 14122 25707 14156 25741
rect 14122 25635 14156 25669
rect 14122 25563 14156 25597
rect 14122 25491 14156 25525
rect 14122 25419 14156 25453
rect 14122 25347 14156 25381
rect 14122 25275 14156 25309
rect 14122 25203 14156 25237
rect 14122 25131 14156 25165
rect 14122 25059 14156 25093
rect 14122 24987 14156 25021
rect 14122 24915 14156 24949
rect 14122 24843 14156 24877
rect 14122 24771 14156 24805
rect 14122 24699 14156 24733
rect 14122 24627 14156 24661
rect 14122 24555 14156 24589
rect 14122 24483 14156 24517
rect 14122 24411 14156 24445
rect 14122 24339 14156 24373
rect 14122 24267 14156 24301
rect 14122 24195 14156 24229
rect 14122 24123 14156 24157
rect 14122 24051 14156 24085
rect 14122 23979 14156 24013
rect 14122 23907 14156 23941
rect 14122 23835 14156 23869
rect 14122 23763 14156 23797
rect 14122 23691 14156 23725
rect 14122 23619 14156 23653
rect 14122 23547 14156 23581
rect 14122 23475 14156 23509
rect 14122 23403 14156 23437
rect 14122 23331 14156 23365
rect 14122 23259 14156 23293
rect 14122 23187 14156 23221
rect 14122 23115 14156 23149
rect 14122 23043 14156 23077
rect 14122 22971 14156 23005
rect 14122 22899 14156 22933
rect 14122 22827 14156 22861
rect 14122 22755 14156 22789
rect 14122 22683 14156 22717
rect 14122 22611 14156 22645
rect 14122 22539 14156 22573
rect 14122 22467 14156 22501
rect 14122 22395 14156 22429
rect 14122 22323 14156 22357
rect 14122 22251 14156 22285
rect 14122 22179 14156 22213
rect 14122 22107 14156 22141
rect 14122 22035 14156 22069
rect 14122 21963 14156 21997
rect 14122 21891 14156 21925
rect 14122 21819 14156 21853
rect 14122 21747 14156 21781
rect 14122 21675 14156 21709
rect 14122 21603 14156 21637
rect 14122 21531 14156 21565
rect 14122 21459 14156 21493
rect 14122 21387 14156 21421
rect 14122 21315 14156 21349
rect 14122 21243 14156 21277
rect 14122 21171 14156 21205
rect 14122 21099 14156 21133
rect 14122 21027 14156 21061
rect 14122 20955 14156 20989
rect 14122 20883 14156 20917
rect 14122 20811 14156 20845
rect 14122 20739 14156 20773
rect 14122 20667 14156 20701
rect 14122 20595 14156 20629
rect 14122 20523 14156 20557
rect 14122 20451 14156 20485
rect 14122 20379 14156 20413
rect 14122 20307 14156 20341
rect 14122 20235 14156 20269
rect 14122 20163 14156 20197
rect 14122 20091 14156 20125
rect 14122 20019 14156 20053
rect 14122 19947 14156 19981
rect 14122 19875 14156 19909
rect 14122 19803 14156 19837
rect 14122 19731 14156 19765
rect 14122 19659 14156 19693
rect 14122 19587 14156 19621
rect 14122 19515 14156 19549
rect 14122 19443 14156 19477
rect 14122 19371 14156 19405
rect 14122 19299 14156 19333
rect 14122 19227 14156 19261
rect 14122 19155 14156 19189
rect 14122 19083 14156 19117
rect 14122 19011 14156 19045
rect 14122 18939 14156 18973
rect 14122 18867 14156 18901
rect 14122 18795 14156 18829
rect 14122 18723 14156 18757
rect 14122 18651 14156 18685
rect 14122 18579 14156 18613
rect 14122 18507 14156 18541
rect 14122 18435 14156 18469
rect 14122 18363 14156 18397
rect 14122 18291 14156 18325
rect 14122 18219 14156 18253
rect 14122 18147 14156 18181
rect 14122 18075 14156 18109
rect 14122 18003 14156 18037
rect 14122 17931 14156 17965
rect 14122 17859 14156 17893
rect 14122 17787 14156 17821
rect 14122 17715 14156 17749
rect 14122 17643 14156 17677
rect 14122 17571 14156 17605
rect 14122 17499 14156 17533
rect 14122 17427 14156 17461
rect 14122 17355 14156 17389
rect 14122 17283 14156 17317
rect 14122 17211 14156 17245
rect 14122 17139 14156 17173
rect 14122 17067 14156 17101
rect 14122 16995 14156 17029
rect 14122 16923 14156 16957
rect 14122 16851 14156 16885
rect 14122 16779 14156 16813
rect 14122 16707 14156 16741
rect 14122 16635 14156 16669
rect 14122 16563 14156 16597
rect 14122 16491 14156 16525
rect 14122 16419 14156 16453
rect 14122 16347 14156 16381
rect 14122 16275 14156 16309
rect 14122 16203 14156 16237
rect 14122 16131 14156 16165
rect 14122 16059 14156 16093
rect 14122 15987 14156 16021
rect 14122 15915 14156 15949
rect 14122 15843 14156 15877
rect 14122 15771 14156 15805
rect 14122 15699 14156 15733
rect 14122 15627 14156 15661
rect 14122 15555 14156 15589
rect 14122 15483 14156 15517
rect 14122 15411 14156 15445
rect 14122 15339 14156 15373
rect 14122 15267 14156 15301
rect 807 15130 841 15164
rect 807 15058 841 15092
rect 14122 15195 14156 15229
rect 14122 15123 14156 15157
rect 14122 15051 14156 15085
rect 891 14908 925 14942
rect 963 14908 997 14942
rect 1035 14908 1069 14942
rect 1107 14908 1141 14942
rect 1179 14908 1213 14942
rect 1251 14908 1285 14942
rect 1323 14908 1357 14942
rect 1395 14908 1429 14942
rect 1467 14908 1501 14942
rect 1539 14908 1573 14942
rect 1611 14908 1645 14942
rect 1683 14908 1717 14942
rect 1755 14908 1789 14942
rect 1827 14908 1861 14942
rect 1899 14908 1933 14942
rect 1971 14908 2005 14942
rect 2043 14908 2077 14942
rect 2115 14908 2149 14942
rect 2187 14908 2221 14942
rect 2259 14908 2293 14942
rect 2331 14908 2365 14942
rect 2403 14908 2437 14942
rect 2475 14908 2509 14942
rect 2547 14908 2581 14942
rect 2619 14908 2653 14942
rect 2691 14908 2725 14942
rect 2763 14908 2797 14942
rect 2835 14908 2869 14942
rect 2907 14908 2941 14942
rect 2979 14908 3013 14942
rect 3051 14908 3085 14942
rect 3123 14908 3157 14942
rect 3195 14908 3229 14942
rect 3267 14908 3301 14942
rect 3339 14908 3373 14942
rect 3411 14908 3445 14942
rect 3483 14908 3517 14942
rect 3555 14908 3589 14942
rect 3627 14908 3661 14942
rect 3699 14908 3733 14942
rect 3771 14908 3805 14942
rect 3843 14908 3877 14942
rect 3915 14908 3949 14942
rect 3987 14908 4021 14942
rect 4059 14908 4093 14942
rect 4131 14908 4165 14942
rect 4203 14908 4237 14942
rect 4275 14908 4309 14942
rect 4347 14908 4381 14942
rect 4419 14908 4453 14942
rect 4491 14908 4525 14942
rect 4563 14908 4597 14942
rect 4635 14908 4669 14942
rect 4707 14908 4741 14942
rect 4779 14908 4813 14942
rect 4851 14908 4885 14942
rect 4923 14908 4957 14942
rect 4995 14908 5029 14942
rect 5067 14908 5101 14942
rect 5139 14908 5173 14942
rect 5211 14908 5245 14942
rect 5283 14908 5317 14942
rect 5355 14908 5389 14942
rect 5427 14908 5461 14942
rect 5499 14908 5533 14942
rect 5571 14908 5605 14942
rect 5643 14908 5677 14942
rect 5715 14908 5749 14942
rect 5787 14908 5821 14942
rect 5859 14908 5893 14942
rect 5931 14908 5965 14942
rect 6003 14908 6037 14942
rect 6075 14908 6109 14942
rect 6147 14908 6181 14942
rect 6219 14908 6253 14942
rect 6291 14908 6325 14942
rect 6363 14908 6397 14942
rect 6435 14908 6469 14942
rect 6507 14908 6541 14942
rect 6579 14908 6613 14942
rect 6651 14908 6685 14942
rect 6723 14908 6757 14942
rect 6795 14908 6829 14942
rect 6867 14908 6901 14942
rect 6939 14908 6973 14942
rect 7011 14908 7045 14942
rect 7083 14908 7117 14942
rect 7155 14908 7189 14942
rect 7227 14908 7261 14942
rect 7299 14908 7333 14942
rect 7371 14908 7405 14942
rect 7443 14908 7477 14942
rect 7515 14908 7549 14942
rect 7587 14908 7621 14942
rect 7659 14908 7693 14942
rect 7731 14908 7765 14942
rect 7803 14908 7837 14942
rect 7875 14908 7909 14942
rect 7947 14908 7981 14942
rect 8019 14908 8053 14942
rect 8091 14908 8125 14942
rect 8163 14908 8197 14942
rect 8235 14908 8269 14942
rect 8307 14908 8341 14942
rect 8379 14908 8413 14942
rect 8451 14908 8485 14942
rect 8523 14908 8557 14942
rect 8595 14908 8629 14942
rect 8667 14908 8701 14942
rect 8739 14908 8773 14942
rect 8811 14908 8845 14942
rect 8883 14908 8917 14942
rect 8955 14908 8989 14942
rect 9027 14908 9061 14942
rect 9099 14908 9133 14942
rect 9171 14908 9205 14942
rect 9243 14908 9277 14942
rect 9315 14908 9349 14942
rect 9387 14908 9421 14942
rect 9459 14908 9493 14942
rect 9531 14908 9565 14942
rect 9603 14908 9637 14942
rect 9675 14908 9709 14942
rect 9747 14908 9781 14942
rect 9819 14908 9853 14942
rect 9891 14908 9925 14942
rect 9963 14908 9997 14942
rect 10035 14908 10069 14942
rect 10107 14908 10141 14942
rect 10179 14908 10213 14942
rect 10251 14908 10285 14942
rect 10323 14908 10357 14942
rect 10395 14908 10429 14942
rect 10467 14908 10501 14942
rect 10539 14908 10573 14942
rect 10611 14908 10645 14942
rect 10683 14908 10717 14942
rect 10755 14908 10789 14942
rect 10827 14908 10861 14942
rect 10899 14908 10933 14942
rect 10971 14908 11005 14942
rect 11043 14908 11077 14942
rect 11115 14908 11149 14942
rect 11187 14908 11221 14942
rect 11259 14908 11293 14942
rect 11331 14908 11365 14942
rect 11403 14908 11437 14942
rect 11475 14908 11509 14942
rect 11547 14908 11581 14942
rect 11619 14908 11653 14942
rect 11691 14908 11725 14942
rect 11763 14908 11797 14942
rect 11835 14908 11869 14942
rect 11907 14908 11941 14942
rect 11979 14908 12013 14942
rect 12051 14908 12085 14942
rect 12123 14908 12157 14942
rect 12195 14908 12229 14942
rect 12267 14908 12301 14942
rect 12339 14908 12373 14942
rect 12411 14908 12445 14942
rect 12483 14908 12517 14942
rect 12555 14908 12589 14942
rect 12627 14908 12661 14942
rect 12699 14908 12733 14942
rect 12771 14908 12805 14942
rect 12843 14908 12877 14942
rect 12915 14908 12949 14942
rect 12987 14908 13021 14942
rect 13059 14908 13093 14942
rect 13131 14908 13165 14942
rect 13203 14908 13237 14942
rect 13275 14908 13309 14942
rect 13347 14908 13381 14942
rect 13419 14908 13453 14942
rect 13491 14908 13525 14942
rect 13563 14908 13597 14942
rect 13635 14908 13669 14942
rect 13707 14908 13741 14942
rect 13779 14908 13813 14942
rect 13851 14908 13885 14942
rect 13923 14908 13957 14942
rect 13995 14908 14029 14942
rect 883 14741 902 14774
rect 902 14741 917 14774
rect 955 14741 970 14774
rect 970 14741 989 14774
rect 1027 14741 1038 14774
rect 1038 14741 1061 14774
rect 1099 14741 1106 14774
rect 1106 14741 1133 14774
rect 1171 14741 1174 14774
rect 1174 14741 1205 14774
rect 1243 14741 1276 14774
rect 1276 14741 1277 14774
rect 1315 14741 1344 14774
rect 1344 14741 1349 14774
rect 1387 14741 1412 14774
rect 1412 14741 1421 14774
rect 1459 14741 1480 14774
rect 1480 14741 1493 14774
rect 1531 14741 1548 14774
rect 1548 14741 1565 14774
rect 1603 14741 1616 14774
rect 1616 14741 1637 14774
rect 1675 14741 1684 14774
rect 1684 14741 1709 14774
rect 1747 14741 1752 14774
rect 1752 14741 1781 14774
rect 1819 14741 1820 14774
rect 1820 14741 1853 14774
rect 1891 14741 1922 14774
rect 1922 14741 1925 14774
rect 1963 14741 1990 14774
rect 1990 14741 1997 14774
rect 2035 14741 2058 14774
rect 2058 14741 2069 14774
rect 12883 14741 12904 14774
rect 12904 14741 12917 14774
rect 12955 14741 12972 14774
rect 12972 14741 12989 14774
rect 13027 14741 13040 14774
rect 13040 14741 13061 14774
rect 13099 14741 13108 14774
rect 13108 14741 13133 14774
rect 13171 14741 13176 14774
rect 13176 14741 13205 14774
rect 13243 14741 13244 14774
rect 13244 14741 13277 14774
rect 13315 14741 13346 14774
rect 13346 14741 13349 14774
rect 13387 14741 13414 14774
rect 13414 14741 13421 14774
rect 13459 14741 13482 14774
rect 13482 14741 13493 14774
rect 13531 14741 13550 14774
rect 13550 14741 13565 14774
rect 13603 14741 13618 14774
rect 13618 14741 13637 14774
rect 13675 14741 13686 14774
rect 13686 14741 13709 14774
rect 13747 14741 13754 14774
rect 13754 14741 13781 14774
rect 13819 14741 13822 14774
rect 13822 14741 13853 14774
rect 13891 14741 13924 14774
rect 13924 14741 13925 14774
rect 13963 14741 13992 14774
rect 13992 14741 13997 14774
rect 14035 14741 14060 14774
rect 14060 14741 14069 14774
rect 883 14740 917 14741
rect 955 14740 989 14741
rect 1027 14740 1061 14741
rect 1099 14740 1133 14741
rect 1171 14740 1205 14741
rect 1243 14740 1277 14741
rect 1315 14740 1349 14741
rect 1387 14740 1421 14741
rect 1459 14740 1493 14741
rect 1531 14740 1565 14741
rect 1603 14740 1637 14741
rect 1675 14740 1709 14741
rect 1747 14740 1781 14741
rect 1819 14740 1853 14741
rect 1891 14740 1925 14741
rect 1963 14740 1997 14741
rect 2035 14740 2069 14741
rect 12883 14740 12917 14741
rect 12955 14740 12989 14741
rect 13027 14740 13061 14741
rect 13099 14740 13133 14741
rect 13171 14740 13205 14741
rect 13243 14740 13277 14741
rect 13315 14740 13349 14741
rect 13387 14740 13421 14741
rect 13459 14740 13493 14741
rect 13531 14740 13565 14741
rect 13603 14740 13637 14741
rect 13675 14740 13709 14741
rect 13747 14740 13781 14741
rect 13819 14740 13853 14741
rect 13891 14740 13925 14741
rect 13963 14740 13997 14741
rect 14035 14740 14069 14741
rect 14614 36192 14641 36206
rect 14641 36192 14648 36206
rect 14614 36172 14648 36192
rect 14614 36124 14641 36134
rect 14641 36124 14648 36134
rect 14614 36100 14648 36124
rect 14614 36056 14641 36062
rect 14641 36056 14648 36062
rect 14614 36028 14648 36056
rect 14614 35988 14641 35990
rect 14641 35988 14648 35990
rect 14614 35956 14648 35988
rect 14614 35886 14648 35918
rect 14614 35884 14641 35886
rect 14641 35884 14648 35886
rect 14614 35818 14648 35846
rect 14614 35812 14641 35818
rect 14641 35812 14648 35818
rect 14614 35750 14648 35774
rect 14614 35740 14641 35750
rect 14641 35740 14648 35750
rect 14614 35682 14648 35702
rect 14614 35668 14641 35682
rect 14641 35668 14648 35682
rect 14614 35614 14648 35630
rect 14614 35596 14641 35614
rect 14641 35596 14648 35614
rect 14614 35546 14648 35558
rect 14614 35524 14641 35546
rect 14641 35524 14648 35546
rect 14614 35478 14648 35486
rect 14614 35452 14641 35478
rect 14641 35452 14648 35478
rect 14614 35410 14648 35414
rect 14614 35380 14641 35410
rect 14641 35380 14648 35410
rect 14614 35308 14641 35342
rect 14641 35308 14648 35342
rect 14614 35240 14641 35270
rect 14641 35240 14648 35270
rect 14614 35236 14648 35240
rect 14614 35172 14641 35198
rect 14641 35172 14648 35198
rect 14614 35164 14648 35172
rect 14614 35104 14641 35126
rect 14641 35104 14648 35126
rect 14614 35092 14648 35104
rect 14614 35036 14641 35054
rect 14641 35036 14648 35054
rect 14614 35020 14648 35036
rect 14614 34968 14641 34982
rect 14641 34968 14648 34982
rect 14614 34948 14648 34968
rect 14614 34900 14641 34910
rect 14641 34900 14648 34910
rect 14614 34876 14648 34900
rect 14614 34832 14641 34838
rect 14641 34832 14648 34838
rect 14614 34804 14648 34832
rect 14614 34764 14641 34766
rect 14641 34764 14648 34766
rect 14614 34732 14648 34764
rect 14614 34662 14648 34694
rect 14614 34660 14641 34662
rect 14641 34660 14648 34662
rect 14614 34594 14648 34622
rect 14614 34588 14641 34594
rect 14641 34588 14648 34594
rect 14614 34526 14648 34550
rect 14614 34516 14641 34526
rect 14641 34516 14648 34526
rect 14614 34458 14648 34478
rect 14614 34444 14641 34458
rect 14641 34444 14648 34458
rect 14614 34390 14648 34406
rect 14614 34372 14641 34390
rect 14641 34372 14648 34390
rect 14614 34322 14648 34334
rect 14614 34300 14641 34322
rect 14641 34300 14648 34322
rect 14614 34254 14648 34262
rect 14614 34228 14641 34254
rect 14641 34228 14648 34254
rect 14614 34186 14648 34190
rect 14614 34156 14641 34186
rect 14641 34156 14648 34186
rect 14614 34084 14641 34118
rect 14641 34084 14648 34118
rect 14614 34016 14641 34046
rect 14641 34016 14648 34046
rect 14614 34012 14648 34016
rect 14614 33948 14641 33974
rect 14641 33948 14648 33974
rect 14614 33940 14648 33948
rect 14614 33880 14641 33902
rect 14641 33880 14648 33902
rect 14614 33868 14648 33880
rect 14614 33812 14641 33830
rect 14641 33812 14648 33830
rect 14614 33796 14648 33812
rect 14614 33744 14641 33758
rect 14641 33744 14648 33758
rect 14614 33724 14648 33744
rect 14614 33676 14641 33686
rect 14641 33676 14648 33686
rect 14614 33652 14648 33676
rect 14614 33608 14641 33614
rect 14641 33608 14648 33614
rect 14614 33580 14648 33608
rect 14614 33540 14641 33542
rect 14641 33540 14648 33542
rect 14614 33508 14648 33540
rect 14614 33438 14648 33470
rect 14614 33436 14641 33438
rect 14641 33436 14648 33438
rect 14614 33370 14648 33398
rect 14614 33364 14641 33370
rect 14641 33364 14648 33370
rect 14614 33302 14648 33326
rect 14614 33292 14641 33302
rect 14641 33292 14648 33302
rect 14614 33234 14648 33254
rect 14614 33220 14641 33234
rect 14641 33220 14648 33234
rect 14614 33166 14648 33182
rect 14614 33148 14641 33166
rect 14641 33148 14648 33166
rect 14614 33098 14648 33110
rect 14614 33076 14641 33098
rect 14641 33076 14648 33098
rect 14614 33030 14648 33038
rect 14614 33004 14641 33030
rect 14641 33004 14648 33030
rect 14614 32962 14648 32966
rect 14614 32932 14641 32962
rect 14641 32932 14648 32962
rect 14614 32860 14641 32894
rect 14641 32860 14648 32894
rect 14614 32792 14641 32822
rect 14641 32792 14648 32822
rect 14614 32788 14648 32792
rect 14614 32724 14641 32750
rect 14641 32724 14648 32750
rect 14614 32716 14648 32724
rect 14614 32656 14641 32678
rect 14641 32656 14648 32678
rect 14614 32644 14648 32656
rect 14614 32588 14641 32606
rect 14641 32588 14648 32606
rect 14614 32572 14648 32588
rect 14614 32520 14641 32534
rect 14641 32520 14648 32534
rect 14614 32500 14648 32520
rect 14614 32452 14641 32462
rect 14641 32452 14648 32462
rect 14614 32428 14648 32452
rect 14614 32384 14641 32390
rect 14641 32384 14648 32390
rect 14614 32356 14648 32384
rect 14614 32316 14641 32318
rect 14641 32316 14648 32318
rect 14614 32284 14648 32316
rect 14614 32214 14648 32246
rect 14614 32212 14641 32214
rect 14641 32212 14648 32214
rect 14614 32146 14648 32174
rect 14614 32140 14641 32146
rect 14641 32140 14648 32146
rect 14614 32078 14648 32102
rect 14614 32068 14641 32078
rect 14641 32068 14648 32078
rect 14614 32010 14648 32030
rect 14614 31996 14641 32010
rect 14641 31996 14648 32010
rect 14614 31942 14648 31958
rect 14614 31924 14641 31942
rect 14641 31924 14648 31942
rect 14614 31874 14648 31886
rect 14614 31852 14641 31874
rect 14641 31852 14648 31874
rect 14614 31806 14648 31814
rect 14614 31780 14641 31806
rect 14641 31780 14648 31806
rect 14614 31738 14648 31742
rect 14614 31708 14641 31738
rect 14641 31708 14648 31738
rect 14614 31636 14641 31670
rect 14641 31636 14648 31670
rect 14614 31568 14641 31598
rect 14641 31568 14648 31598
rect 14614 31564 14648 31568
rect 14614 31500 14641 31526
rect 14641 31500 14648 31526
rect 14614 31492 14648 31500
rect 14614 31432 14641 31454
rect 14641 31432 14648 31454
rect 14614 31420 14648 31432
rect 14614 31364 14641 31382
rect 14641 31364 14648 31382
rect 14614 31348 14648 31364
rect 14614 31296 14641 31310
rect 14641 31296 14648 31310
rect 14614 31276 14648 31296
rect 14614 31228 14641 31238
rect 14641 31228 14648 31238
rect 14614 31204 14648 31228
rect 14614 31160 14641 31166
rect 14641 31160 14648 31166
rect 14614 31132 14648 31160
rect 14614 31092 14641 31094
rect 14641 31092 14648 31094
rect 14614 31060 14648 31092
rect 14614 30990 14648 31022
rect 14614 30988 14641 30990
rect 14641 30988 14648 30990
rect 14614 30922 14648 30950
rect 14614 30916 14641 30922
rect 14641 30916 14648 30922
rect 14614 30854 14648 30878
rect 14614 30844 14641 30854
rect 14641 30844 14648 30854
rect 14614 30786 14648 30806
rect 14614 30772 14641 30786
rect 14641 30772 14648 30786
rect 14614 30718 14648 30734
rect 14614 30700 14641 30718
rect 14641 30700 14648 30718
rect 14614 30650 14648 30662
rect 14614 30628 14641 30650
rect 14641 30628 14648 30650
rect 14614 30582 14648 30590
rect 14614 30556 14641 30582
rect 14641 30556 14648 30582
rect 14614 30514 14648 30518
rect 14614 30484 14641 30514
rect 14641 30484 14648 30514
rect 14614 30412 14641 30446
rect 14641 30412 14648 30446
rect 14614 30344 14641 30374
rect 14641 30344 14648 30374
rect 14614 30340 14648 30344
rect 14614 30276 14641 30302
rect 14641 30276 14648 30302
rect 14614 30268 14648 30276
rect 14614 30208 14641 30230
rect 14641 30208 14648 30230
rect 14614 30196 14648 30208
rect 14614 30140 14641 30158
rect 14641 30140 14648 30158
rect 14614 30124 14648 30140
rect 14614 30072 14641 30086
rect 14641 30072 14648 30086
rect 14614 30052 14648 30072
rect 14614 30004 14641 30014
rect 14641 30004 14648 30014
rect 14614 29980 14648 30004
rect 14614 29936 14641 29942
rect 14641 29936 14648 29942
rect 14614 29908 14648 29936
rect 14614 29868 14641 29870
rect 14641 29868 14648 29870
rect 14614 29836 14648 29868
rect 14614 29766 14648 29798
rect 14614 29764 14641 29766
rect 14641 29764 14648 29766
rect 14614 29698 14648 29726
rect 14614 29692 14641 29698
rect 14641 29692 14648 29698
rect 14614 29630 14648 29654
rect 14614 29620 14641 29630
rect 14641 29620 14648 29630
rect 14614 29562 14648 29582
rect 14614 29548 14641 29562
rect 14641 29548 14648 29562
rect 14614 29494 14648 29510
rect 14614 29476 14641 29494
rect 14641 29476 14648 29494
rect 14614 29426 14648 29438
rect 14614 29404 14641 29426
rect 14641 29404 14648 29426
rect 14614 29358 14648 29366
rect 14614 29332 14641 29358
rect 14641 29332 14648 29358
rect 14614 29290 14648 29294
rect 14614 29260 14641 29290
rect 14641 29260 14648 29290
rect 14614 29188 14641 29222
rect 14641 29188 14648 29222
rect 14614 29120 14641 29150
rect 14641 29120 14648 29150
rect 14614 29116 14648 29120
rect 14614 29052 14641 29078
rect 14641 29052 14648 29078
rect 14614 29044 14648 29052
rect 14614 28984 14641 29006
rect 14641 28984 14648 29006
rect 14614 28972 14648 28984
rect 14614 28916 14641 28934
rect 14641 28916 14648 28934
rect 14614 28900 14648 28916
rect 14614 28848 14641 28862
rect 14641 28848 14648 28862
rect 14614 28828 14648 28848
rect 14614 28780 14641 28790
rect 14641 28780 14648 28790
rect 14614 28756 14648 28780
rect 14614 28712 14641 28718
rect 14641 28712 14648 28718
rect 14614 28684 14648 28712
rect 14614 28644 14641 28646
rect 14641 28644 14648 28646
rect 14614 28612 14648 28644
rect 14614 28542 14648 28574
rect 14614 28540 14641 28542
rect 14641 28540 14648 28542
rect 14614 28474 14648 28502
rect 14614 28468 14641 28474
rect 14641 28468 14648 28474
rect 14614 28406 14648 28430
rect 14614 28396 14641 28406
rect 14641 28396 14648 28406
rect 14614 28338 14648 28358
rect 14614 28324 14641 28338
rect 14641 28324 14648 28338
rect 14614 28270 14648 28286
rect 14614 28252 14641 28270
rect 14641 28252 14648 28270
rect 14614 28202 14648 28214
rect 14614 28180 14641 28202
rect 14641 28180 14648 28202
rect 14614 28134 14648 28142
rect 14614 28108 14641 28134
rect 14641 28108 14648 28134
rect 14614 28066 14648 28070
rect 14614 28036 14641 28066
rect 14641 28036 14648 28066
rect 14614 27964 14641 27998
rect 14641 27964 14648 27998
rect 14614 27896 14641 27926
rect 14641 27896 14648 27926
rect 14614 27892 14648 27896
rect 14614 27828 14641 27854
rect 14641 27828 14648 27854
rect 14614 27820 14648 27828
rect 14614 27760 14641 27782
rect 14641 27760 14648 27782
rect 14614 27748 14648 27760
rect 14614 27692 14641 27710
rect 14641 27692 14648 27710
rect 14614 27676 14648 27692
rect 14614 27624 14641 27638
rect 14641 27624 14648 27638
rect 14614 27604 14648 27624
rect 14614 27556 14641 27566
rect 14641 27556 14648 27566
rect 14614 27532 14648 27556
rect 14614 27488 14641 27494
rect 14641 27488 14648 27494
rect 14614 27460 14648 27488
rect 14614 27420 14641 27422
rect 14641 27420 14648 27422
rect 14614 27388 14648 27420
rect 14614 27318 14648 27350
rect 14614 27316 14641 27318
rect 14641 27316 14648 27318
rect 14614 27250 14648 27278
rect 14614 27244 14641 27250
rect 14641 27244 14648 27250
rect 14614 27182 14648 27206
rect 14614 27172 14641 27182
rect 14641 27172 14648 27182
rect 14614 27114 14648 27134
rect 14614 27100 14641 27114
rect 14641 27100 14648 27114
rect 14614 27046 14648 27062
rect 14614 27028 14641 27046
rect 14641 27028 14648 27046
rect 14614 26978 14648 26990
rect 14614 26956 14641 26978
rect 14641 26956 14648 26978
rect 14614 26910 14648 26918
rect 14614 26884 14641 26910
rect 14641 26884 14648 26910
rect 14614 26842 14648 26846
rect 14614 26812 14641 26842
rect 14641 26812 14648 26842
rect 14614 26740 14641 26774
rect 14641 26740 14648 26774
rect 14614 26672 14641 26702
rect 14641 26672 14648 26702
rect 14614 26668 14648 26672
rect 14614 26604 14641 26630
rect 14641 26604 14648 26630
rect 14614 26596 14648 26604
rect 14614 26536 14641 26558
rect 14641 26536 14648 26558
rect 14614 26524 14648 26536
rect 14614 26468 14641 26486
rect 14641 26468 14648 26486
rect 14614 26452 14648 26468
rect 14614 26400 14641 26414
rect 14641 26400 14648 26414
rect 14614 26380 14648 26400
rect 14614 26332 14641 26342
rect 14641 26332 14648 26342
rect 14614 26308 14648 26332
rect 14614 26264 14641 26270
rect 14641 26264 14648 26270
rect 14614 26236 14648 26264
rect 14614 26196 14641 26198
rect 14641 26196 14648 26198
rect 14614 26164 14648 26196
rect 14614 26094 14648 26126
rect 14614 26092 14641 26094
rect 14641 26092 14648 26094
rect 14614 26026 14648 26054
rect 14614 26020 14641 26026
rect 14641 26020 14648 26026
rect 14614 25958 14648 25982
rect 14614 25948 14641 25958
rect 14641 25948 14648 25958
rect 14614 25890 14648 25910
rect 14614 25876 14641 25890
rect 14641 25876 14648 25890
rect 14614 25822 14648 25838
rect 14614 25804 14641 25822
rect 14641 25804 14648 25822
rect 14614 25754 14648 25766
rect 14614 25732 14641 25754
rect 14641 25732 14648 25754
rect 14614 25686 14648 25694
rect 14614 25660 14641 25686
rect 14641 25660 14648 25686
rect 14614 25618 14648 25622
rect 14614 25588 14641 25618
rect 14641 25588 14648 25618
rect 14614 25516 14641 25550
rect 14641 25516 14648 25550
rect 14614 25448 14641 25478
rect 14641 25448 14648 25478
rect 14614 25444 14648 25448
rect 14614 25380 14641 25406
rect 14641 25380 14648 25406
rect 14614 25372 14648 25380
rect 14614 25312 14641 25334
rect 14641 25312 14648 25334
rect 14614 25300 14648 25312
rect 14614 25244 14641 25262
rect 14641 25244 14648 25262
rect 14614 25228 14648 25244
rect 14614 25176 14641 25190
rect 14641 25176 14648 25190
rect 14614 25156 14648 25176
rect 14614 25108 14641 25118
rect 14641 25108 14648 25118
rect 14614 25084 14648 25108
rect 14614 25040 14641 25046
rect 14641 25040 14648 25046
rect 14614 25012 14648 25040
rect 14614 24972 14641 24974
rect 14641 24972 14648 24974
rect 14614 24940 14648 24972
rect 14614 24870 14648 24902
rect 14614 24868 14641 24870
rect 14641 24868 14648 24870
rect 14614 24802 14648 24830
rect 14614 24796 14641 24802
rect 14641 24796 14648 24802
rect 14614 24734 14648 24758
rect 14614 24724 14641 24734
rect 14641 24724 14648 24734
rect 14614 24666 14648 24686
rect 14614 24652 14641 24666
rect 14641 24652 14648 24666
rect 14614 24598 14648 24614
rect 14614 24580 14641 24598
rect 14641 24580 14648 24598
rect 14614 24530 14648 24542
rect 14614 24508 14641 24530
rect 14641 24508 14648 24530
rect 14614 24462 14648 24470
rect 14614 24436 14641 24462
rect 14641 24436 14648 24462
rect 14614 24394 14648 24398
rect 14614 24364 14641 24394
rect 14641 24364 14648 24394
rect 14614 24292 14641 24326
rect 14641 24292 14648 24326
rect 14614 24224 14641 24254
rect 14641 24224 14648 24254
rect 14614 24220 14648 24224
rect 14614 24156 14641 24182
rect 14641 24156 14648 24182
rect 14614 24148 14648 24156
rect 14614 24088 14641 24110
rect 14641 24088 14648 24110
rect 14614 24076 14648 24088
rect 14614 24020 14641 24038
rect 14641 24020 14648 24038
rect 14614 24004 14648 24020
rect 14614 23952 14641 23966
rect 14641 23952 14648 23966
rect 14614 23932 14648 23952
rect 14614 23884 14641 23894
rect 14641 23884 14648 23894
rect 14614 23860 14648 23884
rect 14614 23816 14641 23822
rect 14641 23816 14648 23822
rect 14614 23788 14648 23816
rect 14614 23748 14641 23750
rect 14641 23748 14648 23750
rect 14614 23716 14648 23748
rect 14614 23646 14648 23678
rect 14614 23644 14641 23646
rect 14641 23644 14648 23646
rect 14614 23578 14648 23606
rect 14614 23572 14641 23578
rect 14641 23572 14648 23578
rect 14614 23510 14648 23534
rect 14614 23500 14641 23510
rect 14641 23500 14648 23510
rect 14614 23442 14648 23462
rect 14614 23428 14641 23442
rect 14641 23428 14648 23442
rect 14614 23374 14648 23390
rect 14614 23356 14641 23374
rect 14641 23356 14648 23374
rect 14614 23306 14648 23318
rect 14614 23284 14641 23306
rect 14641 23284 14648 23306
rect 14614 23238 14648 23246
rect 14614 23212 14641 23238
rect 14641 23212 14648 23238
rect 14614 23170 14648 23174
rect 14614 23140 14641 23170
rect 14641 23140 14648 23170
rect 14614 23068 14641 23102
rect 14641 23068 14648 23102
rect 14614 23000 14641 23030
rect 14641 23000 14648 23030
rect 14614 22996 14648 23000
rect 14614 22932 14641 22958
rect 14641 22932 14648 22958
rect 14614 22924 14648 22932
rect 14614 22864 14641 22886
rect 14641 22864 14648 22886
rect 14614 22852 14648 22864
rect 14614 22796 14641 22814
rect 14641 22796 14648 22814
rect 14614 22780 14648 22796
rect 14614 22728 14641 22742
rect 14641 22728 14648 22742
rect 14614 22708 14648 22728
rect 14614 22660 14641 22670
rect 14641 22660 14648 22670
rect 14614 22636 14648 22660
rect 14614 22592 14641 22598
rect 14641 22592 14648 22598
rect 14614 22564 14648 22592
rect 14614 22524 14641 22526
rect 14641 22524 14648 22526
rect 14614 22492 14648 22524
rect 14614 22422 14648 22454
rect 14614 22420 14641 22422
rect 14641 22420 14648 22422
rect 14614 22354 14648 22382
rect 14614 22348 14641 22354
rect 14641 22348 14648 22354
rect 14614 22286 14648 22310
rect 14614 22276 14641 22286
rect 14641 22276 14648 22286
rect 14614 22218 14648 22238
rect 14614 22204 14641 22218
rect 14641 22204 14648 22218
rect 14614 22150 14648 22166
rect 14614 22132 14641 22150
rect 14641 22132 14648 22150
rect 14614 22082 14648 22094
rect 14614 22060 14641 22082
rect 14641 22060 14648 22082
rect 14614 22014 14648 22022
rect 14614 21988 14641 22014
rect 14641 21988 14648 22014
rect 14614 21946 14648 21950
rect 14614 21916 14641 21946
rect 14641 21916 14648 21946
rect 14614 21844 14641 21878
rect 14641 21844 14648 21878
rect 14614 21776 14641 21806
rect 14641 21776 14648 21806
rect 14614 21772 14648 21776
rect 14614 21708 14641 21734
rect 14641 21708 14648 21734
rect 14614 21700 14648 21708
rect 14614 21640 14641 21662
rect 14641 21640 14648 21662
rect 14614 21628 14648 21640
rect 14614 21572 14641 21590
rect 14641 21572 14648 21590
rect 14614 21556 14648 21572
rect 14614 21504 14641 21518
rect 14641 21504 14648 21518
rect 14614 21484 14648 21504
rect 14614 21436 14641 21446
rect 14641 21436 14648 21446
rect 14614 21412 14648 21436
rect 14614 21368 14641 21374
rect 14641 21368 14648 21374
rect 14614 21340 14648 21368
rect 14614 21300 14641 21302
rect 14641 21300 14648 21302
rect 14614 21268 14648 21300
rect 14614 21198 14648 21230
rect 14614 21196 14641 21198
rect 14641 21196 14648 21198
rect 14614 21130 14648 21158
rect 14614 21124 14641 21130
rect 14641 21124 14648 21130
rect 14614 21062 14648 21086
rect 14614 21052 14641 21062
rect 14641 21052 14648 21062
rect 14614 20994 14648 21014
rect 14614 20980 14641 20994
rect 14641 20980 14648 20994
rect 14614 20926 14648 20942
rect 14614 20908 14641 20926
rect 14641 20908 14648 20926
rect 14614 20858 14648 20870
rect 14614 20836 14641 20858
rect 14641 20836 14648 20858
rect 14614 20790 14648 20798
rect 14614 20764 14641 20790
rect 14641 20764 14648 20790
rect 14614 20722 14648 20726
rect 14614 20692 14641 20722
rect 14641 20692 14648 20722
rect 14614 20620 14641 20654
rect 14641 20620 14648 20654
rect 14614 20552 14641 20582
rect 14641 20552 14648 20582
rect 14614 20548 14648 20552
rect 14614 20484 14641 20510
rect 14641 20484 14648 20510
rect 14614 20476 14648 20484
rect 14614 20416 14641 20438
rect 14641 20416 14648 20438
rect 14614 20404 14648 20416
rect 14614 20348 14641 20366
rect 14641 20348 14648 20366
rect 14614 20332 14648 20348
rect 14614 20280 14641 20294
rect 14641 20280 14648 20294
rect 14614 20260 14648 20280
rect 14614 20212 14641 20222
rect 14641 20212 14648 20222
rect 14614 20188 14648 20212
rect 14614 20144 14641 20150
rect 14641 20144 14648 20150
rect 14614 20116 14648 20144
rect 14614 20076 14641 20078
rect 14641 20076 14648 20078
rect 14614 20044 14648 20076
rect 14614 19974 14648 20006
rect 14614 19972 14641 19974
rect 14641 19972 14648 19974
rect 14614 19906 14648 19934
rect 14614 19900 14641 19906
rect 14641 19900 14648 19906
rect 14614 19838 14648 19862
rect 14614 19828 14641 19838
rect 14641 19828 14648 19838
rect 14614 19770 14648 19790
rect 14614 19756 14641 19770
rect 14641 19756 14648 19770
rect 14614 19702 14648 19718
rect 14614 19684 14641 19702
rect 14641 19684 14648 19702
rect 14614 19634 14648 19646
rect 14614 19612 14641 19634
rect 14641 19612 14648 19634
rect 14614 19566 14648 19574
rect 14614 19540 14641 19566
rect 14641 19540 14648 19566
rect 14614 19498 14648 19502
rect 14614 19468 14641 19498
rect 14641 19468 14648 19498
rect 14614 19396 14641 19430
rect 14641 19396 14648 19430
rect 14614 19328 14641 19358
rect 14641 19328 14648 19358
rect 14614 19324 14648 19328
rect 14614 19260 14641 19286
rect 14641 19260 14648 19286
rect 14614 19252 14648 19260
rect 14614 19192 14641 19214
rect 14641 19192 14648 19214
rect 14614 19180 14648 19192
rect 14614 19124 14641 19142
rect 14641 19124 14648 19142
rect 14614 19108 14648 19124
rect 14614 19056 14641 19070
rect 14641 19056 14648 19070
rect 14614 19036 14648 19056
rect 14614 18988 14641 18998
rect 14641 18988 14648 18998
rect 14614 18964 14648 18988
rect 14614 18920 14641 18926
rect 14641 18920 14648 18926
rect 14614 18892 14648 18920
rect 14614 18852 14641 18854
rect 14641 18852 14648 18854
rect 14614 18820 14648 18852
rect 14614 18750 14648 18782
rect 14614 18748 14641 18750
rect 14641 18748 14648 18750
rect 14614 18682 14648 18710
rect 14614 18676 14641 18682
rect 14641 18676 14648 18682
rect 14614 18614 14648 18638
rect 14614 18604 14641 18614
rect 14641 18604 14648 18614
rect 14614 18546 14648 18566
rect 14614 18532 14641 18546
rect 14641 18532 14648 18546
rect 14614 18478 14648 18494
rect 14614 18460 14641 18478
rect 14641 18460 14648 18478
rect 14614 18410 14648 18422
rect 14614 18388 14641 18410
rect 14641 18388 14648 18410
rect 14614 18342 14648 18350
rect 14614 18316 14641 18342
rect 14641 18316 14648 18342
rect 14614 18274 14648 18278
rect 14614 18244 14641 18274
rect 14641 18244 14648 18274
rect 14614 18172 14641 18206
rect 14641 18172 14648 18206
rect 14614 18104 14641 18134
rect 14641 18104 14648 18134
rect 14614 18100 14648 18104
rect 14614 18036 14641 18062
rect 14641 18036 14648 18062
rect 14614 18028 14648 18036
rect 14614 17968 14641 17990
rect 14641 17968 14648 17990
rect 14614 17956 14648 17968
rect 14614 17900 14641 17918
rect 14641 17900 14648 17918
rect 14614 17884 14648 17900
rect 14614 17832 14641 17846
rect 14641 17832 14648 17846
rect 14614 17812 14648 17832
rect 14614 17764 14641 17774
rect 14641 17764 14648 17774
rect 14614 17740 14648 17764
rect 14614 17696 14641 17702
rect 14641 17696 14648 17702
rect 14614 17668 14648 17696
rect 14614 17628 14641 17630
rect 14641 17628 14648 17630
rect 14614 17596 14648 17628
rect 14614 17526 14648 17558
rect 14614 17524 14641 17526
rect 14641 17524 14648 17526
rect 14614 17458 14648 17486
rect 14614 17452 14641 17458
rect 14641 17452 14648 17458
rect 14614 17390 14648 17414
rect 14614 17380 14641 17390
rect 14641 17380 14648 17390
rect 14614 17322 14648 17342
rect 14614 17308 14641 17322
rect 14641 17308 14648 17322
rect 14614 17254 14648 17270
rect 14614 17236 14641 17254
rect 14641 17236 14648 17254
rect 14614 17186 14648 17198
rect 14614 17164 14641 17186
rect 14641 17164 14648 17186
rect 14614 17118 14648 17126
rect 14614 17092 14641 17118
rect 14641 17092 14648 17118
rect 14614 17050 14648 17054
rect 14614 17020 14641 17050
rect 14641 17020 14648 17050
rect 14614 16948 14641 16982
rect 14641 16948 14648 16982
rect 14614 16880 14641 16910
rect 14641 16880 14648 16910
rect 14614 16876 14648 16880
rect 14614 16812 14641 16838
rect 14641 16812 14648 16838
rect 14614 16804 14648 16812
rect 14614 16744 14641 16766
rect 14641 16744 14648 16766
rect 14614 16732 14648 16744
rect 14614 16676 14641 16694
rect 14641 16676 14648 16694
rect 14614 16660 14648 16676
rect 14614 16608 14641 16622
rect 14641 16608 14648 16622
rect 14614 16588 14648 16608
rect 14614 16540 14641 16550
rect 14641 16540 14648 16550
rect 14614 16516 14648 16540
rect 14614 16472 14641 16478
rect 14641 16472 14648 16478
rect 14614 16444 14648 16472
rect 14614 16404 14641 16406
rect 14641 16404 14648 16406
rect 14614 16372 14648 16404
rect 14614 16302 14648 16334
rect 14614 16300 14641 16302
rect 14641 16300 14648 16302
rect 14614 16234 14648 16262
rect 14614 16228 14641 16234
rect 14641 16228 14648 16234
rect 14614 16166 14648 16190
rect 14614 16156 14641 16166
rect 14641 16156 14648 16166
rect 14614 16098 14648 16118
rect 14614 16084 14641 16098
rect 14641 16084 14648 16098
rect 14614 16030 14648 16046
rect 14614 16012 14641 16030
rect 14641 16012 14648 16030
rect 14614 15962 14648 15974
rect 14614 15940 14641 15962
rect 14641 15940 14648 15962
rect 14614 15894 14648 15902
rect 14614 15868 14641 15894
rect 14641 15868 14648 15894
rect 14614 15826 14648 15830
rect 14614 15796 14641 15826
rect 14641 15796 14648 15826
rect 14614 15724 14641 15758
rect 14641 15724 14648 15758
rect 14614 15656 14641 15686
rect 14641 15656 14648 15686
rect 14614 15652 14648 15656
rect 14614 15588 14641 15614
rect 14641 15588 14648 15614
rect 14614 15580 14648 15588
rect 14614 15520 14641 15542
rect 14641 15520 14648 15542
rect 14614 15508 14648 15520
rect 14614 15452 14641 15470
rect 14641 15452 14648 15470
rect 14614 15436 14648 15452
rect 14614 15384 14641 15398
rect 14641 15384 14648 15398
rect 14614 15364 14648 15384
rect 14614 15316 14641 15326
rect 14641 15316 14648 15326
rect 14614 15292 14648 15316
rect 14614 15248 14641 15254
rect 14641 15248 14648 15254
rect 14614 15220 14648 15248
rect 14614 15180 14641 15182
rect 14641 15180 14648 15182
rect 14614 15148 14648 15180
rect 14614 15078 14648 15110
rect 14614 15076 14641 15078
rect 14641 15076 14648 15078
rect 14614 15010 14648 15038
rect 14614 15004 14641 15010
rect 14641 15004 14648 15010
rect 14614 14942 14648 14966
rect 14614 14932 14641 14942
rect 14641 14932 14648 14942
rect 14614 14874 14648 14894
rect 14614 14860 14641 14874
rect 14641 14860 14648 14874
rect 14614 14806 14648 14822
rect 14614 14788 14641 14806
rect 14641 14788 14648 14806
rect 14614 14738 14648 14750
rect 320 14664 354 14681
rect 320 14647 346 14664
rect 346 14647 354 14664
rect 14614 14716 14641 14738
rect 14641 14716 14648 14738
rect 14614 14670 14648 14678
rect 14614 14644 14641 14670
rect 14641 14644 14648 14670
rect 320 14418 354 14452
rect 610 14451 644 14452
rect 2311 14451 2345 14452
rect 2383 14451 2417 14452
rect 2455 14451 2489 14452
rect 2527 14451 2561 14452
rect 2599 14451 2633 14452
rect 2671 14451 2705 14452
rect 2743 14451 2777 14452
rect 2815 14451 2849 14452
rect 2887 14451 2921 14452
rect 2959 14451 2993 14452
rect 3031 14451 3065 14452
rect 3103 14451 3137 14452
rect 3175 14451 3209 14452
rect 3247 14451 3281 14452
rect 3319 14451 3353 14452
rect 3391 14451 3425 14452
rect 3463 14451 3497 14452
rect 3535 14451 3569 14452
rect 3607 14451 3641 14452
rect 3679 14451 3713 14452
rect 3751 14451 3785 14452
rect 3823 14451 3857 14452
rect 3895 14451 3929 14452
rect 3967 14451 4001 14452
rect 4039 14451 4073 14452
rect 4111 14451 4145 14452
rect 4183 14451 4217 14452
rect 4255 14451 4289 14452
rect 4327 14451 4361 14452
rect 4399 14451 4433 14452
rect 4471 14451 4505 14452
rect 4543 14451 4577 14452
rect 4615 14451 4649 14452
rect 4687 14451 4721 14452
rect 4759 14451 4793 14452
rect 4831 14451 4865 14452
rect 4903 14451 4937 14452
rect 4975 14451 5009 14452
rect 5047 14451 5081 14452
rect 5119 14451 5153 14452
rect 5191 14451 5225 14452
rect 5263 14451 5297 14452
rect 5335 14451 5369 14452
rect 5407 14451 5441 14452
rect 5479 14451 5513 14452
rect 5551 14451 5585 14452
rect 5623 14451 5657 14452
rect 5695 14451 5729 14452
rect 5767 14451 5801 14452
rect 5839 14451 5873 14452
rect 5911 14451 5945 14452
rect 5983 14451 6017 14452
rect 6055 14451 6089 14452
rect 6127 14451 6161 14452
rect 6199 14451 6233 14452
rect 6271 14451 6305 14452
rect 6343 14451 6377 14452
rect 6415 14451 6449 14452
rect 6487 14451 6521 14452
rect 6559 14451 6593 14452
rect 6631 14451 6665 14452
rect 6703 14451 6737 14452
rect 6775 14451 6809 14452
rect 6847 14451 6881 14452
rect 6919 14451 6953 14452
rect 6991 14451 7025 14452
rect 7063 14451 7097 14452
rect 7135 14451 7169 14452
rect 7207 14451 7241 14452
rect 7279 14451 7313 14452
rect 7351 14451 7385 14452
rect 7423 14451 7457 14452
rect 7495 14451 7529 14452
rect 7567 14451 7601 14452
rect 7639 14451 7673 14452
rect 7711 14451 7745 14452
rect 7783 14451 7817 14452
rect 7855 14451 7889 14452
rect 7927 14451 7961 14452
rect 7999 14451 8033 14452
rect 8071 14451 8105 14452
rect 8143 14451 8177 14452
rect 8215 14451 8249 14452
rect 8287 14451 8321 14452
rect 8359 14451 8393 14452
rect 8431 14451 8465 14452
rect 8503 14451 8537 14452
rect 8575 14451 8609 14452
rect 8647 14451 8681 14452
rect 8719 14451 8753 14452
rect 8791 14451 8825 14452
rect 8863 14451 8897 14452
rect 8935 14451 8969 14452
rect 9007 14451 9041 14452
rect 9079 14451 9113 14452
rect 9151 14451 9185 14452
rect 9223 14451 9257 14452
rect 9295 14451 9329 14452
rect 9367 14451 9401 14452
rect 9439 14451 9473 14452
rect 9511 14451 9545 14452
rect 9583 14451 9617 14452
rect 9655 14451 9689 14452
rect 9727 14451 9761 14452
rect 9799 14451 9833 14452
rect 9871 14451 9905 14452
rect 9943 14451 9977 14452
rect 10015 14451 10049 14452
rect 10087 14451 10121 14452
rect 10159 14451 10193 14452
rect 10231 14451 10265 14452
rect 10303 14451 10337 14452
rect 10375 14451 10409 14452
rect 10447 14451 10481 14452
rect 10519 14451 10553 14452
rect 10591 14451 10625 14452
rect 10663 14451 10697 14452
rect 10735 14451 10769 14452
rect 10807 14451 10841 14452
rect 10879 14451 10913 14452
rect 10951 14451 10985 14452
rect 11023 14451 11057 14452
rect 11095 14451 11129 14452
rect 11167 14451 11201 14452
rect 11239 14451 11273 14452
rect 11311 14451 11345 14452
rect 11383 14451 11417 14452
rect 11455 14451 11489 14452
rect 11527 14451 11561 14452
rect 11599 14451 11633 14452
rect 11671 14451 11705 14452
rect 11743 14451 11777 14452
rect 11815 14451 11849 14452
rect 11887 14451 11921 14452
rect 11959 14451 11993 14452
rect 12031 14451 12065 14452
rect 12103 14451 12137 14452
rect 12175 14451 12209 14452
rect 12247 14451 12281 14452
rect 12319 14451 12353 14452
rect 12391 14451 12425 14452
rect 12463 14451 12497 14452
rect 12535 14451 12569 14452
rect 12607 14451 12641 14452
rect 610 14418 612 14451
rect 612 14418 644 14451
rect 2311 14418 2312 14451
rect 2312 14418 2345 14451
rect 2383 14418 2414 14451
rect 2414 14418 2417 14451
rect 2455 14418 2482 14451
rect 2482 14418 2489 14451
rect 2527 14418 2550 14451
rect 2550 14418 2561 14451
rect 2599 14418 2618 14451
rect 2618 14418 2633 14451
rect 2671 14418 2686 14451
rect 2686 14418 2705 14451
rect 2743 14418 2754 14451
rect 2754 14418 2777 14451
rect 2815 14418 2822 14451
rect 2822 14418 2849 14451
rect 2887 14418 2890 14451
rect 2890 14418 2921 14451
rect 2959 14418 2992 14451
rect 2992 14418 2993 14451
rect 3031 14418 3060 14451
rect 3060 14418 3065 14451
rect 3103 14418 3128 14451
rect 3128 14418 3137 14451
rect 3175 14418 3196 14451
rect 3196 14418 3209 14451
rect 3247 14418 3264 14451
rect 3264 14418 3281 14451
rect 3319 14418 3332 14451
rect 3332 14418 3353 14451
rect 3391 14418 3400 14451
rect 3400 14418 3425 14451
rect 3463 14418 3468 14451
rect 3468 14418 3497 14451
rect 3535 14418 3536 14451
rect 3536 14418 3569 14451
rect 3607 14418 3638 14451
rect 3638 14418 3641 14451
rect 3679 14418 3706 14451
rect 3706 14418 3713 14451
rect 3751 14418 3774 14451
rect 3774 14418 3785 14451
rect 3823 14418 3842 14451
rect 3842 14418 3857 14451
rect 3895 14418 3910 14451
rect 3910 14418 3929 14451
rect 3967 14418 3978 14451
rect 3978 14418 4001 14451
rect 4039 14418 4046 14451
rect 4046 14418 4073 14451
rect 4111 14418 4114 14451
rect 4114 14418 4145 14451
rect 4183 14418 4216 14451
rect 4216 14418 4217 14451
rect 4255 14418 4284 14451
rect 4284 14418 4289 14451
rect 4327 14418 4352 14451
rect 4352 14418 4361 14451
rect 4399 14418 4420 14451
rect 4420 14418 4433 14451
rect 4471 14418 4488 14451
rect 4488 14418 4505 14451
rect 4543 14418 4556 14451
rect 4556 14418 4577 14451
rect 4615 14418 4624 14451
rect 4624 14418 4649 14451
rect 4687 14418 4692 14451
rect 4692 14418 4721 14451
rect 4759 14418 4760 14451
rect 4760 14418 4793 14451
rect 4831 14418 4862 14451
rect 4862 14418 4865 14451
rect 4903 14418 4930 14451
rect 4930 14418 4937 14451
rect 4975 14418 4998 14451
rect 4998 14418 5009 14451
rect 5047 14418 5066 14451
rect 5066 14418 5081 14451
rect 5119 14418 5134 14451
rect 5134 14418 5153 14451
rect 5191 14418 5202 14451
rect 5202 14418 5225 14451
rect 5263 14418 5270 14451
rect 5270 14418 5297 14451
rect 5335 14418 5338 14451
rect 5338 14418 5369 14451
rect 5407 14418 5440 14451
rect 5440 14418 5441 14451
rect 5479 14418 5508 14451
rect 5508 14418 5513 14451
rect 5551 14418 5576 14451
rect 5576 14418 5585 14451
rect 5623 14418 5644 14451
rect 5644 14418 5657 14451
rect 5695 14418 5712 14451
rect 5712 14418 5729 14451
rect 5767 14418 5780 14451
rect 5780 14418 5801 14451
rect 5839 14418 5848 14451
rect 5848 14418 5873 14451
rect 5911 14418 5916 14451
rect 5916 14418 5945 14451
rect 5983 14418 5984 14451
rect 5984 14418 6017 14451
rect 6055 14418 6086 14451
rect 6086 14418 6089 14451
rect 6127 14418 6154 14451
rect 6154 14418 6161 14451
rect 6199 14418 6222 14451
rect 6222 14418 6233 14451
rect 6271 14418 6290 14451
rect 6290 14418 6305 14451
rect 6343 14418 6358 14451
rect 6358 14418 6377 14451
rect 6415 14418 6426 14451
rect 6426 14418 6449 14451
rect 6487 14418 6494 14451
rect 6494 14418 6521 14451
rect 6559 14418 6562 14451
rect 6562 14418 6593 14451
rect 6631 14418 6664 14451
rect 6664 14418 6665 14451
rect 6703 14418 6732 14451
rect 6732 14418 6737 14451
rect 6775 14418 6800 14451
rect 6800 14418 6809 14451
rect 6847 14418 6868 14451
rect 6868 14418 6881 14451
rect 6919 14418 6936 14451
rect 6936 14418 6953 14451
rect 6991 14418 7004 14451
rect 7004 14418 7025 14451
rect 7063 14418 7072 14451
rect 7072 14418 7097 14451
rect 7135 14418 7140 14451
rect 7140 14418 7169 14451
rect 7207 14418 7208 14451
rect 7208 14418 7241 14451
rect 7279 14418 7310 14451
rect 7310 14418 7313 14451
rect 7351 14418 7378 14451
rect 7378 14418 7385 14451
rect 7423 14418 7446 14451
rect 7446 14418 7457 14451
rect 7495 14418 7514 14451
rect 7514 14418 7529 14451
rect 7567 14418 7582 14451
rect 7582 14418 7601 14451
rect 7639 14418 7650 14451
rect 7650 14418 7673 14451
rect 7711 14418 7718 14451
rect 7718 14418 7745 14451
rect 7783 14418 7786 14451
rect 7786 14418 7817 14451
rect 7855 14418 7888 14451
rect 7888 14418 7889 14451
rect 7927 14418 7956 14451
rect 7956 14418 7961 14451
rect 7999 14418 8024 14451
rect 8024 14418 8033 14451
rect 8071 14418 8092 14451
rect 8092 14418 8105 14451
rect 8143 14418 8160 14451
rect 8160 14418 8177 14451
rect 8215 14418 8228 14451
rect 8228 14418 8249 14451
rect 8287 14418 8296 14451
rect 8296 14418 8321 14451
rect 8359 14418 8364 14451
rect 8364 14418 8393 14451
rect 8431 14418 8432 14451
rect 8432 14418 8465 14451
rect 8503 14418 8534 14451
rect 8534 14418 8537 14451
rect 8575 14418 8602 14451
rect 8602 14418 8609 14451
rect 8647 14418 8670 14451
rect 8670 14418 8681 14451
rect 8719 14418 8738 14451
rect 8738 14418 8753 14451
rect 8791 14418 8806 14451
rect 8806 14418 8825 14451
rect 8863 14418 8874 14451
rect 8874 14418 8897 14451
rect 8935 14418 8942 14451
rect 8942 14418 8969 14451
rect 9007 14418 9010 14451
rect 9010 14418 9041 14451
rect 9079 14418 9112 14451
rect 9112 14418 9113 14451
rect 9151 14418 9180 14451
rect 9180 14418 9185 14451
rect 9223 14418 9248 14451
rect 9248 14418 9257 14451
rect 9295 14418 9316 14451
rect 9316 14418 9329 14451
rect 9367 14418 9384 14451
rect 9384 14418 9401 14451
rect 9439 14418 9452 14451
rect 9452 14418 9473 14451
rect 9511 14418 9520 14451
rect 9520 14418 9545 14451
rect 9583 14418 9588 14451
rect 9588 14418 9617 14451
rect 9655 14418 9656 14451
rect 9656 14418 9689 14451
rect 9727 14418 9758 14451
rect 9758 14418 9761 14451
rect 9799 14418 9826 14451
rect 9826 14418 9833 14451
rect 9871 14418 9894 14451
rect 9894 14418 9905 14451
rect 9943 14418 9962 14451
rect 9962 14418 9977 14451
rect 10015 14418 10030 14451
rect 10030 14418 10049 14451
rect 10087 14418 10098 14451
rect 10098 14418 10121 14451
rect 10159 14418 10166 14451
rect 10166 14418 10193 14451
rect 10231 14418 10234 14451
rect 10234 14418 10265 14451
rect 10303 14418 10336 14451
rect 10336 14418 10337 14451
rect 10375 14418 10404 14451
rect 10404 14418 10409 14451
rect 10447 14418 10472 14451
rect 10472 14418 10481 14451
rect 10519 14418 10540 14451
rect 10540 14418 10553 14451
rect 10591 14418 10608 14451
rect 10608 14418 10625 14451
rect 10663 14418 10676 14451
rect 10676 14418 10697 14451
rect 10735 14418 10744 14451
rect 10744 14418 10769 14451
rect 10807 14418 10812 14451
rect 10812 14418 10841 14451
rect 10879 14418 10880 14451
rect 10880 14418 10913 14451
rect 10951 14418 10982 14451
rect 10982 14418 10985 14451
rect 11023 14418 11050 14451
rect 11050 14418 11057 14451
rect 11095 14418 11118 14451
rect 11118 14418 11129 14451
rect 11167 14418 11186 14451
rect 11186 14418 11201 14451
rect 11239 14418 11254 14451
rect 11254 14418 11273 14451
rect 11311 14418 11322 14451
rect 11322 14418 11345 14451
rect 11383 14418 11390 14451
rect 11390 14418 11417 14451
rect 11455 14418 11458 14451
rect 11458 14418 11489 14451
rect 11527 14418 11560 14451
rect 11560 14418 11561 14451
rect 11599 14418 11628 14451
rect 11628 14418 11633 14451
rect 11671 14418 11696 14451
rect 11696 14418 11705 14451
rect 11743 14418 11764 14451
rect 11764 14418 11777 14451
rect 11815 14418 11832 14451
rect 11832 14418 11849 14451
rect 11887 14418 11900 14451
rect 11900 14418 11921 14451
rect 11959 14418 11968 14451
rect 11968 14418 11993 14451
rect 12031 14418 12036 14451
rect 12036 14418 12065 14451
rect 12103 14418 12104 14451
rect 12104 14418 12137 14451
rect 12175 14418 12206 14451
rect 12206 14418 12209 14451
rect 12247 14418 12274 14451
rect 12274 14418 12281 14451
rect 12319 14418 12342 14451
rect 12342 14418 12353 14451
rect 12391 14418 12410 14451
rect 12410 14418 12425 14451
rect 12463 14418 12478 14451
rect 12478 14418 12497 14451
rect 12535 14418 12546 14451
rect 12546 14418 12569 14451
rect 12607 14418 12614 14451
rect 12614 14418 12641 14451
rect 14314 14418 14348 14452
rect 14614 14418 14648 14452
<< metal1 >>
rect 885 37211 2234 37258
rect 885 36574 957 37211
rect 245 36534 957 36574
rect 245 36500 320 36534
rect 354 36500 957 36534
rect 245 36498 957 36500
rect 2161 36574 2234 37211
rect 12752 37208 14101 37262
rect 12752 36574 12821 37208
rect 2161 36498 12821 36574
rect 14025 36574 14101 37208
rect 14025 36533 14724 36574
rect 14025 36499 14614 36533
rect 14648 36499 14724 36533
rect 14025 36498 14724 36499
rect 245 36464 556 36498
rect 590 36464 628 36498
rect 662 36464 700 36498
rect 734 36464 772 36498
rect 806 36464 844 36498
rect 878 36464 916 36498
rect 950 36464 957 36498
rect 2174 36464 2212 36498
rect 2246 36464 2284 36498
rect 2318 36464 2356 36498
rect 2390 36464 2428 36498
rect 2462 36464 2500 36498
rect 2534 36464 2572 36498
rect 2606 36464 2644 36498
rect 2678 36464 2716 36498
rect 2750 36464 2788 36498
rect 2822 36464 2860 36498
rect 2894 36464 2932 36498
rect 2966 36464 3004 36498
rect 3038 36464 3076 36498
rect 3110 36464 3148 36498
rect 3182 36464 3220 36498
rect 3254 36464 3292 36498
rect 3326 36464 3364 36498
rect 3398 36464 3436 36498
rect 3470 36464 3508 36498
rect 3542 36464 3580 36498
rect 3614 36464 3652 36498
rect 3686 36464 3724 36498
rect 3758 36464 3796 36498
rect 3830 36464 3868 36498
rect 3902 36464 3940 36498
rect 3974 36464 4012 36498
rect 4046 36464 4084 36498
rect 4118 36464 4156 36498
rect 4190 36464 4228 36498
rect 4262 36464 4300 36498
rect 4334 36464 4372 36498
rect 4406 36464 4444 36498
rect 4478 36464 4516 36498
rect 4550 36464 4588 36498
rect 4622 36464 4660 36498
rect 4694 36464 4732 36498
rect 4766 36464 4804 36498
rect 4838 36464 4876 36498
rect 4910 36464 4948 36498
rect 4982 36464 5020 36498
rect 5054 36464 5092 36498
rect 5126 36464 5164 36498
rect 5198 36464 5236 36498
rect 5270 36464 5308 36498
rect 5342 36464 5380 36498
rect 5414 36464 5452 36498
rect 5486 36464 5524 36498
rect 5558 36464 5596 36498
rect 5630 36464 5668 36498
rect 5702 36464 5740 36498
rect 5774 36464 5812 36498
rect 5846 36464 5884 36498
rect 5918 36464 5956 36498
rect 5990 36464 6028 36498
rect 6062 36464 6100 36498
rect 6134 36464 6172 36498
rect 6206 36464 6244 36498
rect 6278 36464 6316 36498
rect 6350 36464 6388 36498
rect 6422 36464 6460 36498
rect 6494 36464 6532 36498
rect 6566 36464 6604 36498
rect 6638 36464 6676 36498
rect 6710 36464 6748 36498
rect 6782 36464 6820 36498
rect 6854 36464 6892 36498
rect 6926 36464 6964 36498
rect 6998 36464 7036 36498
rect 7070 36464 7108 36498
rect 7142 36464 7180 36498
rect 7214 36464 7252 36498
rect 7286 36464 7324 36498
rect 7358 36464 7396 36498
rect 7430 36464 7468 36498
rect 7502 36464 7540 36498
rect 7574 36464 7612 36498
rect 7646 36464 7684 36498
rect 7718 36464 7756 36498
rect 7790 36464 7828 36498
rect 7862 36464 7900 36498
rect 7934 36464 7972 36498
rect 8006 36464 8044 36498
rect 8078 36464 8116 36498
rect 8150 36464 8188 36498
rect 8222 36464 8260 36498
rect 8294 36464 8332 36498
rect 8366 36464 8404 36498
rect 8438 36464 8476 36498
rect 8510 36464 8548 36498
rect 8582 36464 8620 36498
rect 8654 36464 8692 36498
rect 8726 36464 8764 36498
rect 8798 36464 8836 36498
rect 8870 36464 8908 36498
rect 8942 36464 8980 36498
rect 9014 36464 9052 36498
rect 9086 36464 9124 36498
rect 9158 36464 9196 36498
rect 9230 36464 9268 36498
rect 9302 36464 9340 36498
rect 9374 36464 9412 36498
rect 9446 36464 9484 36498
rect 9518 36464 9556 36498
rect 9590 36464 9628 36498
rect 9662 36464 9700 36498
rect 9734 36464 9772 36498
rect 9806 36464 9844 36498
rect 9878 36464 9916 36498
rect 9950 36464 9988 36498
rect 10022 36464 10060 36498
rect 10094 36464 10132 36498
rect 10166 36464 10204 36498
rect 10238 36464 10276 36498
rect 10310 36464 10348 36498
rect 10382 36464 10420 36498
rect 10454 36464 10492 36498
rect 10526 36464 10564 36498
rect 10598 36464 10636 36498
rect 10670 36464 10708 36498
rect 10742 36464 10780 36498
rect 10814 36464 10852 36498
rect 10886 36464 10924 36498
rect 10958 36464 10996 36498
rect 11030 36464 11068 36498
rect 11102 36464 11140 36498
rect 11174 36464 11212 36498
rect 11246 36464 11284 36498
rect 11318 36464 11356 36498
rect 11390 36464 11428 36498
rect 11462 36464 11500 36498
rect 11534 36464 11572 36498
rect 11606 36464 11644 36498
rect 11678 36464 11716 36498
rect 11750 36464 11788 36498
rect 11822 36464 11860 36498
rect 11894 36464 11932 36498
rect 11966 36464 12004 36498
rect 12038 36464 12076 36498
rect 12110 36464 12148 36498
rect 12182 36464 12220 36498
rect 12254 36464 12292 36498
rect 12326 36464 12364 36498
rect 12398 36464 12436 36498
rect 12470 36464 12508 36498
rect 12542 36464 12580 36498
rect 12614 36464 12652 36498
rect 12686 36464 12724 36498
rect 12758 36464 12796 36498
rect 14054 36464 14092 36498
rect 14126 36464 14164 36498
rect 14198 36464 14236 36498
rect 14270 36464 14308 36498
rect 14342 36464 14380 36498
rect 14414 36464 14724 36498
rect 245 36462 957 36464
rect 245 36428 320 36462
rect 354 36455 957 36462
rect 2161 36455 12821 36464
rect 354 36452 12821 36455
rect 14025 36461 14724 36464
rect 14025 36452 14614 36461
rect 354 36428 14614 36452
rect 245 36427 14614 36428
rect 14648 36427 14724 36461
rect 245 36389 14724 36427
rect 245 36281 430 36389
rect 245 36247 320 36281
rect 354 36247 430 36281
rect 245 36209 430 36247
rect 245 36175 320 36209
rect 354 36175 430 36209
rect 245 36137 430 36175
rect 245 36103 320 36137
rect 354 36103 430 36137
rect 245 36065 430 36103
rect 245 36031 320 36065
rect 354 36031 430 36065
rect 14539 36278 14724 36389
rect 14539 36244 14614 36278
rect 14648 36244 14724 36278
rect 14539 36206 14724 36244
rect 14539 36172 14614 36206
rect 14648 36172 14724 36206
rect 14539 36134 14724 36172
rect 14539 36100 14614 36134
rect 14648 36100 14724 36134
rect 14539 36062 14724 36100
rect 245 35993 430 36031
tri 832 36028 857 36053 se
rect 857 36028 14119 36053
tri 14119 36028 14144 36053 sw
rect 14539 36028 14614 36062
rect 14648 36028 14724 36062
tri 823 36019 832 36028 se
rect 832 36019 14144 36028
tri 807 36003 823 36019 se
rect 823 36003 14144 36019
rect 245 35959 320 35993
rect 354 35959 430 35993
tri 773 35969 807 36003 se
rect 807 35969 1009 36003
rect 1043 35969 1081 36003
rect 1115 35969 1153 36003
rect 1187 35969 1225 36003
rect 1259 35969 1297 36003
rect 1331 35969 1369 36003
rect 1403 35969 1441 36003
rect 1475 35969 1513 36003
rect 1547 35969 1585 36003
rect 1619 35969 1657 36003
rect 1691 35969 1729 36003
rect 1763 35969 1801 36003
rect 1835 35969 1873 36003
rect 1907 35969 1945 36003
rect 1979 35969 2017 36003
rect 2051 35969 2089 36003
rect 2123 35969 2161 36003
rect 2195 35969 2233 36003
rect 2267 35969 2305 36003
rect 2339 35969 2377 36003
rect 2411 35969 2449 36003
rect 2483 35969 2521 36003
rect 2555 35969 2593 36003
rect 2627 35969 2665 36003
rect 2699 35969 2737 36003
rect 2771 35969 2809 36003
rect 2843 35969 2881 36003
rect 2915 35969 2953 36003
rect 2987 35969 3025 36003
rect 3059 35969 3097 36003
rect 3131 35969 3169 36003
rect 3203 35969 3241 36003
rect 3275 35969 3313 36003
rect 3347 35969 3385 36003
rect 3419 35969 3457 36003
rect 3491 35969 3529 36003
rect 3563 35969 3601 36003
rect 3635 35969 3673 36003
rect 3707 35969 3745 36003
rect 3779 35969 3817 36003
rect 3851 35969 3889 36003
rect 3923 35969 3961 36003
rect 3995 35969 4033 36003
rect 4067 35969 4105 36003
rect 4139 35969 4177 36003
rect 4211 35969 4249 36003
rect 4283 35969 4321 36003
rect 4355 35969 4393 36003
rect 4427 35969 4465 36003
rect 4499 35969 4537 36003
rect 4571 35969 4609 36003
rect 4643 35969 4681 36003
rect 4715 35969 4753 36003
rect 4787 35969 4825 36003
rect 4859 35969 4897 36003
rect 4931 35969 4969 36003
rect 5003 35969 5041 36003
rect 5075 35969 5113 36003
rect 5147 35969 5185 36003
rect 5219 35969 5257 36003
rect 5291 35969 5329 36003
rect 5363 35969 5401 36003
rect 5435 35969 5473 36003
rect 5507 35969 5545 36003
rect 5579 35969 5617 36003
rect 5651 35969 5689 36003
rect 5723 35969 5761 36003
rect 5795 35969 5833 36003
rect 5867 35969 5905 36003
rect 5939 35969 5977 36003
rect 6011 35969 6049 36003
rect 6083 35969 6121 36003
rect 6155 35969 6193 36003
rect 6227 35969 6265 36003
rect 6299 35969 6337 36003
rect 6371 35969 6409 36003
rect 6443 35969 6481 36003
rect 6515 35969 6553 36003
rect 6587 35969 6625 36003
rect 6659 35969 6697 36003
rect 6731 35969 6769 36003
rect 6803 35969 6841 36003
rect 6875 35969 6913 36003
rect 6947 35969 6985 36003
rect 7019 35969 7057 36003
rect 7091 35969 7129 36003
rect 7163 35969 7201 36003
rect 7235 35969 7273 36003
rect 7307 35969 7345 36003
rect 7379 35969 7417 36003
rect 7451 35969 7489 36003
rect 7523 35969 7561 36003
rect 7595 35969 7633 36003
rect 7667 35969 7705 36003
rect 7739 35969 7777 36003
rect 7811 35969 7849 36003
rect 7883 35969 7921 36003
rect 7955 35969 7993 36003
rect 8027 35969 8065 36003
rect 8099 35969 8137 36003
rect 8171 35969 8209 36003
rect 8243 35969 8281 36003
rect 8315 35969 8353 36003
rect 8387 35969 8425 36003
rect 8459 35969 8497 36003
rect 8531 35969 8569 36003
rect 8603 35969 8641 36003
rect 8675 35969 8713 36003
rect 8747 35969 8785 36003
rect 8819 35969 8857 36003
rect 8891 35969 8929 36003
rect 8963 35969 9001 36003
rect 9035 35969 9073 36003
rect 9107 35969 9145 36003
rect 9179 35969 9217 36003
rect 9251 35969 9289 36003
rect 9323 35969 9361 36003
rect 9395 35969 9433 36003
rect 9467 35969 9505 36003
rect 9539 35969 9577 36003
rect 9611 35969 9649 36003
rect 9683 35969 9721 36003
rect 9755 35969 9793 36003
rect 9827 35969 9865 36003
rect 9899 35969 9937 36003
rect 9971 35969 10009 36003
rect 10043 35969 10081 36003
rect 10115 35969 10153 36003
rect 10187 35969 10225 36003
rect 10259 35969 10297 36003
rect 10331 35969 10369 36003
rect 10403 35969 10441 36003
rect 10475 35969 10513 36003
rect 10547 35969 10585 36003
rect 10619 35969 10657 36003
rect 10691 35969 10729 36003
rect 10763 35969 10801 36003
rect 10835 35969 10873 36003
rect 10907 35969 10945 36003
rect 10979 35969 11017 36003
rect 11051 35969 11089 36003
rect 11123 35969 11161 36003
rect 11195 35969 11233 36003
rect 11267 35969 11305 36003
rect 11339 35969 11377 36003
rect 11411 35969 11449 36003
rect 11483 35969 11521 36003
rect 11555 35969 11593 36003
rect 11627 35969 11665 36003
rect 11699 35969 11737 36003
rect 11771 35969 11809 36003
rect 11843 35969 11881 36003
rect 11915 35969 11953 36003
rect 11987 35969 12025 36003
rect 12059 35969 12097 36003
rect 12131 35969 12169 36003
rect 12203 35969 12241 36003
rect 12275 35969 12313 36003
rect 12347 35969 12385 36003
rect 12419 35969 12457 36003
rect 12491 35969 12529 36003
rect 12563 35969 12601 36003
rect 12635 35969 12673 36003
rect 12707 35969 12745 36003
rect 12779 35969 12817 36003
rect 12851 35969 12889 36003
rect 12923 35969 12961 36003
rect 12995 35969 13033 36003
rect 13067 35969 13105 36003
rect 13139 35969 13177 36003
rect 13211 35969 13249 36003
rect 13283 35969 13321 36003
rect 13355 35969 13393 36003
rect 13427 35969 13465 36003
rect 13499 35969 13537 36003
rect 13571 35969 13609 36003
rect 13643 35969 13681 36003
rect 13715 35969 13753 36003
rect 13787 35969 13825 36003
rect 13859 35969 13897 36003
rect 13931 35969 13969 36003
rect 14003 35990 14144 36003
tri 14144 35990 14182 36028 sw
rect 14539 35990 14724 36028
rect 14003 35969 14182 35990
rect 245 35921 430 35959
tri 760 35956 773 35969 se
rect 773 35956 14182 35969
tri 14182 35956 14216 35990 sw
rect 14539 35956 14614 35990
rect 14648 35956 14724 35990
rect 245 35887 320 35921
rect 354 35887 430 35921
rect 245 35849 430 35887
rect 245 35815 320 35849
rect 354 35815 430 35849
rect 245 35777 430 35815
rect 245 35743 320 35777
rect 354 35743 430 35777
rect 245 35705 430 35743
rect 245 35671 320 35705
rect 354 35671 430 35705
rect 245 35633 430 35671
rect 245 35599 320 35633
rect 354 35599 430 35633
rect 245 35561 430 35599
rect 245 35527 320 35561
rect 354 35527 430 35561
rect 245 35489 430 35527
rect 245 35455 320 35489
rect 354 35455 430 35489
rect 245 35417 430 35455
rect 245 35383 320 35417
rect 354 35383 430 35417
rect 245 35345 430 35383
rect 245 35311 320 35345
rect 354 35311 430 35345
rect 245 35273 430 35311
rect 245 35239 320 35273
rect 354 35239 430 35273
rect 245 35201 430 35239
rect 245 35167 320 35201
rect 354 35167 430 35201
rect 245 35129 430 35167
rect 245 35095 320 35129
rect 354 35095 430 35129
rect 245 35057 430 35095
rect 245 35023 320 35057
rect 354 35023 430 35057
rect 245 34985 430 35023
rect 245 34951 320 34985
rect 354 34951 430 34985
rect 245 34913 430 34951
rect 245 34879 320 34913
rect 354 34879 430 34913
rect 245 34841 430 34879
rect 245 34807 320 34841
rect 354 34807 430 34841
rect 245 34769 430 34807
rect 245 34735 320 34769
rect 354 34735 430 34769
rect 245 34697 430 34735
rect 245 34663 320 34697
rect 354 34663 430 34697
rect 245 34625 430 34663
rect 245 34591 320 34625
rect 354 34591 430 34625
rect 245 34553 430 34591
rect 245 34519 320 34553
rect 354 34519 430 34553
rect 245 34481 430 34519
rect 245 34447 320 34481
rect 354 34447 430 34481
rect 245 34409 430 34447
rect 245 34375 320 34409
rect 354 34375 430 34409
rect 245 34337 430 34375
rect 245 34303 320 34337
rect 354 34303 430 34337
rect 245 34265 430 34303
rect 245 34231 320 34265
rect 354 34231 430 34265
rect 245 34193 430 34231
rect 245 34159 320 34193
rect 354 34159 430 34193
rect 245 34121 430 34159
rect 245 34087 320 34121
rect 354 34087 430 34121
rect 245 34049 430 34087
rect 245 34015 320 34049
rect 354 34015 430 34049
rect 245 33977 430 34015
rect 245 33943 320 33977
rect 354 33943 430 33977
rect 245 33905 430 33943
rect 245 33871 320 33905
rect 354 33871 430 33905
rect 245 33833 430 33871
rect 245 33799 320 33833
rect 354 33799 430 33833
rect 245 33761 430 33799
rect 245 33727 320 33761
rect 354 33727 430 33761
rect 245 33689 430 33727
rect 245 33655 320 33689
rect 354 33655 430 33689
rect 245 33617 430 33655
rect 245 33583 320 33617
rect 354 33583 430 33617
rect 245 33545 430 33583
rect 245 33511 320 33545
rect 354 33511 430 33545
rect 245 33473 430 33511
rect 245 33439 320 33473
rect 354 33439 430 33473
rect 245 33401 430 33439
rect 245 33367 320 33401
rect 354 33367 430 33401
rect 245 33329 430 33367
rect 245 33295 320 33329
rect 354 33295 430 33329
rect 245 33257 430 33295
rect 245 33223 320 33257
rect 354 33223 430 33257
rect 245 33185 430 33223
rect 245 33151 320 33185
rect 354 33151 430 33185
rect 245 33113 430 33151
rect 245 33079 320 33113
rect 354 33079 430 33113
rect 245 33041 430 33079
rect 245 33007 320 33041
rect 354 33007 430 33041
rect 245 32969 430 33007
rect 245 32935 320 32969
rect 354 32935 430 32969
rect 245 32897 430 32935
rect 245 32863 320 32897
rect 354 32863 430 32897
rect 245 32825 430 32863
rect 245 32791 320 32825
rect 354 32791 430 32825
rect 245 32753 430 32791
rect 245 32719 320 32753
rect 354 32719 430 32753
rect 245 32681 430 32719
rect 245 32647 320 32681
rect 354 32647 430 32681
rect 245 32609 430 32647
rect 245 32575 320 32609
rect 354 32575 430 32609
rect 245 32537 430 32575
rect 245 32503 320 32537
rect 354 32503 430 32537
rect 245 32465 430 32503
rect 245 32431 320 32465
rect 354 32431 430 32465
rect 245 32393 430 32431
rect 245 32359 320 32393
rect 354 32359 430 32393
rect 245 32321 430 32359
rect 245 32287 320 32321
rect 354 32287 430 32321
rect 245 32249 430 32287
rect 245 32215 320 32249
rect 354 32215 430 32249
rect 245 32177 430 32215
rect 245 32143 320 32177
rect 354 32143 430 32177
rect 245 32105 430 32143
rect 245 32071 320 32105
rect 354 32071 430 32105
rect 245 32033 430 32071
rect 245 31999 320 32033
rect 354 31999 430 32033
rect 245 31961 430 31999
rect 245 31927 320 31961
rect 354 31927 430 31961
rect 245 31889 430 31927
rect 245 31855 320 31889
rect 354 31855 430 31889
rect 245 31817 430 31855
rect 245 31783 320 31817
rect 354 31783 430 31817
rect 245 31745 430 31783
rect 245 31711 320 31745
rect 354 31711 430 31745
rect 245 31673 430 31711
rect 245 31639 320 31673
rect 354 31639 430 31673
rect 245 31601 430 31639
rect 245 31567 320 31601
rect 354 31567 430 31601
rect 245 31529 430 31567
rect 245 31495 320 31529
rect 354 31495 430 31529
rect 245 31457 430 31495
rect 245 31423 320 31457
rect 354 31423 430 31457
rect 245 31385 430 31423
rect 245 31351 320 31385
rect 354 31351 430 31385
rect 245 31313 430 31351
rect 245 31279 320 31313
rect 354 31279 430 31313
rect 245 31241 430 31279
rect 245 31207 320 31241
rect 354 31207 430 31241
rect 245 31169 430 31207
rect 245 31135 320 31169
rect 354 31135 430 31169
rect 245 31097 430 31135
rect 245 31063 320 31097
rect 354 31063 430 31097
rect 245 31025 430 31063
rect 245 30991 320 31025
rect 354 30991 430 31025
rect 245 30953 430 30991
rect 245 30919 320 30953
rect 354 30919 430 30953
rect 245 30881 430 30919
rect 245 30847 320 30881
rect 354 30847 430 30881
rect 245 30809 430 30847
rect 245 30775 320 30809
rect 354 30775 430 30809
rect 245 30737 430 30775
rect 245 30703 320 30737
rect 354 30703 430 30737
rect 245 30665 430 30703
rect 245 30631 320 30665
rect 354 30631 430 30665
rect 245 30593 430 30631
rect 245 30559 320 30593
rect 354 30559 430 30593
rect 245 30521 430 30559
rect 245 30487 320 30521
rect 354 30487 430 30521
rect 245 30449 430 30487
rect 245 30415 320 30449
rect 354 30415 430 30449
rect 245 30377 430 30415
rect 245 30343 320 30377
rect 354 30343 430 30377
rect 245 30305 430 30343
rect 245 30271 320 30305
rect 354 30271 430 30305
rect 245 30233 430 30271
rect 245 30199 320 30233
rect 354 30199 430 30233
rect 245 30161 430 30199
rect 245 30127 320 30161
rect 354 30127 430 30161
rect 245 30089 430 30127
rect 245 30055 320 30089
rect 354 30055 430 30089
rect 245 30017 430 30055
rect 245 29983 320 30017
rect 354 29983 430 30017
rect 245 29945 430 29983
rect 245 29911 320 29945
rect 354 29911 430 29945
rect 245 29873 430 29911
rect 245 29839 320 29873
rect 354 29839 430 29873
rect 245 29801 430 29839
rect 245 29767 320 29801
rect 354 29767 430 29801
rect 245 29729 430 29767
rect 245 29695 320 29729
rect 354 29695 430 29729
rect 245 29657 430 29695
rect 245 29623 320 29657
rect 354 29623 430 29657
rect 245 29585 430 29623
rect 245 29551 320 29585
rect 354 29551 430 29585
rect 245 29513 430 29551
rect 245 29479 320 29513
rect 354 29479 430 29513
rect 245 29441 430 29479
rect 245 29407 320 29441
rect 354 29407 430 29441
rect 245 29369 430 29407
rect 245 29335 320 29369
rect 354 29335 430 29369
rect 245 29297 430 29335
rect 245 29263 320 29297
rect 354 29263 430 29297
rect 245 29225 430 29263
rect 245 29191 320 29225
rect 354 29191 430 29225
rect 245 29153 430 29191
rect 245 29119 320 29153
rect 354 29119 430 29153
rect 245 29081 430 29119
rect 245 29047 320 29081
rect 354 29047 430 29081
rect 245 29009 430 29047
rect 245 28975 320 29009
rect 354 28975 430 29009
rect 245 28937 430 28975
rect 245 28903 320 28937
rect 354 28903 430 28937
rect 245 28865 430 28903
rect 245 28831 320 28865
rect 354 28831 430 28865
rect 245 28793 430 28831
rect 245 28759 320 28793
rect 354 28759 430 28793
rect 245 28721 430 28759
rect 245 28687 320 28721
rect 354 28687 430 28721
rect 245 28649 430 28687
rect 245 28615 320 28649
rect 354 28615 430 28649
rect 245 28577 430 28615
rect 245 28543 320 28577
rect 354 28543 430 28577
rect 245 28505 430 28543
rect 245 28471 320 28505
rect 354 28471 430 28505
rect 245 28433 430 28471
rect 245 28399 320 28433
rect 354 28399 430 28433
rect 245 28361 430 28399
rect 245 28327 320 28361
rect 354 28327 430 28361
rect 245 28289 430 28327
rect 245 28255 320 28289
rect 354 28255 430 28289
rect 245 28217 430 28255
rect 245 28183 320 28217
rect 354 28183 430 28217
rect 245 28145 430 28183
rect 245 28111 320 28145
rect 354 28111 430 28145
rect 245 28073 430 28111
rect 245 28039 320 28073
rect 354 28039 430 28073
rect 245 28001 430 28039
rect 245 27967 320 28001
rect 354 27967 430 28001
rect 245 27929 430 27967
rect 245 27895 320 27929
rect 354 27895 430 27929
rect 245 27857 430 27895
rect 245 27823 320 27857
rect 354 27823 430 27857
rect 245 27785 430 27823
rect 245 27751 320 27785
rect 354 27751 430 27785
rect 245 27713 430 27751
rect 245 27679 320 27713
rect 354 27679 430 27713
rect 245 27641 430 27679
rect 245 27607 320 27641
rect 354 27607 430 27641
rect 245 27569 430 27607
rect 245 27535 320 27569
rect 354 27535 430 27569
rect 245 27497 430 27535
rect 245 27463 320 27497
rect 354 27463 430 27497
rect 245 27425 430 27463
rect 245 27391 320 27425
rect 354 27391 430 27425
rect 245 27353 430 27391
rect 245 27319 320 27353
rect 354 27319 430 27353
rect 245 27281 430 27319
rect 245 27247 320 27281
rect 354 27247 430 27281
rect 245 27209 430 27247
rect 245 27175 320 27209
rect 354 27175 430 27209
rect 245 27137 430 27175
rect 245 27103 320 27137
rect 354 27103 430 27137
rect 245 27065 430 27103
rect 245 27031 320 27065
rect 354 27031 430 27065
rect 245 26993 430 27031
rect 245 26959 320 26993
rect 354 26959 430 26993
rect 245 26921 430 26959
rect 245 26887 320 26921
rect 354 26887 430 26921
rect 245 26849 430 26887
rect 245 26815 320 26849
rect 354 26815 430 26849
rect 245 26777 430 26815
rect 245 26743 320 26777
rect 354 26743 430 26777
rect 245 26705 430 26743
rect 245 26671 320 26705
rect 354 26671 430 26705
rect 245 26633 430 26671
rect 245 26599 320 26633
rect 354 26599 430 26633
rect 245 26561 430 26599
rect 245 26527 320 26561
rect 354 26527 430 26561
rect 245 26489 430 26527
rect 245 26455 320 26489
rect 354 26455 430 26489
rect 245 26417 430 26455
rect 245 26383 320 26417
rect 354 26383 430 26417
rect 245 26345 430 26383
rect 245 26311 320 26345
rect 354 26311 430 26345
rect 245 26273 430 26311
rect 245 26239 320 26273
rect 354 26239 430 26273
rect 245 26201 430 26239
rect 245 26167 320 26201
rect 354 26167 430 26201
rect 245 26129 430 26167
rect 245 26095 320 26129
rect 354 26095 430 26129
rect 245 26057 430 26095
rect 245 26023 320 26057
rect 354 26023 430 26057
rect 245 25985 430 26023
rect 245 25951 320 25985
rect 354 25951 430 25985
rect 245 25913 430 25951
rect 245 25879 320 25913
rect 354 25879 430 25913
rect 245 25841 430 25879
rect 245 25807 320 25841
rect 354 25807 430 25841
rect 245 25769 430 25807
rect 245 25735 320 25769
rect 354 25735 430 25769
rect 245 25697 430 25735
rect 245 25663 320 25697
rect 354 25663 430 25697
rect 245 25625 430 25663
rect 245 25591 320 25625
rect 354 25591 430 25625
rect 245 25553 430 25591
rect 245 25519 320 25553
rect 354 25519 430 25553
rect 245 25481 430 25519
rect 245 25447 320 25481
rect 354 25447 430 25481
rect 245 25409 430 25447
rect 245 25375 320 25409
rect 354 25375 430 25409
rect 245 25337 430 25375
rect 245 25303 320 25337
rect 354 25303 430 25337
rect 245 25265 430 25303
rect 245 25231 320 25265
rect 354 25231 430 25265
rect 245 25193 430 25231
rect 245 25159 320 25193
rect 354 25159 430 25193
rect 245 25121 430 25159
rect 245 25087 320 25121
rect 354 25087 430 25121
rect 245 25049 430 25087
rect 245 25015 320 25049
rect 354 25015 430 25049
rect 245 24977 430 25015
rect 245 24943 320 24977
rect 354 24943 430 24977
rect 245 24905 430 24943
rect 245 24871 320 24905
rect 354 24871 430 24905
rect 245 24833 430 24871
rect 245 24799 320 24833
rect 354 24799 430 24833
rect 245 24761 430 24799
rect 245 24727 320 24761
rect 354 24727 430 24761
rect 245 24689 430 24727
rect 245 24655 320 24689
rect 354 24655 430 24689
rect 245 24617 430 24655
rect 245 24583 320 24617
rect 354 24583 430 24617
rect 245 24545 430 24583
rect 245 24511 320 24545
rect 354 24511 430 24545
rect 245 24473 430 24511
rect 245 24439 320 24473
rect 354 24439 430 24473
rect 245 24401 430 24439
rect 245 24367 320 24401
rect 354 24367 430 24401
rect 245 24329 430 24367
rect 245 24295 320 24329
rect 354 24295 430 24329
rect 245 24257 430 24295
rect 245 24223 320 24257
rect 354 24223 430 24257
rect 245 24185 430 24223
rect 245 24151 320 24185
rect 354 24151 430 24185
rect 245 24113 430 24151
rect 245 24079 320 24113
rect 354 24079 430 24113
rect 245 24041 430 24079
rect 245 24007 320 24041
rect 354 24007 430 24041
rect 245 23969 430 24007
rect 245 23935 320 23969
rect 354 23935 430 23969
rect 245 23897 430 23935
rect 245 23863 320 23897
rect 354 23863 430 23897
rect 245 23825 430 23863
rect 245 23791 320 23825
rect 354 23791 430 23825
rect 245 23753 430 23791
rect 245 23719 320 23753
rect 354 23719 430 23753
rect 245 23681 430 23719
rect 245 23647 320 23681
rect 354 23647 430 23681
rect 245 23609 430 23647
rect 245 23575 320 23609
rect 354 23575 430 23609
rect 245 23537 430 23575
rect 245 23503 320 23537
rect 354 23503 430 23537
rect 245 23465 430 23503
rect 245 23431 320 23465
rect 354 23431 430 23465
rect 245 23393 430 23431
rect 245 23359 320 23393
rect 354 23359 430 23393
rect 245 23321 430 23359
rect 245 23287 320 23321
rect 354 23287 430 23321
rect 245 23249 430 23287
rect 245 23215 320 23249
rect 354 23215 430 23249
rect 245 23177 430 23215
rect 245 23143 320 23177
rect 354 23143 430 23177
rect 245 23105 430 23143
rect 245 23071 320 23105
rect 354 23071 430 23105
rect 245 23033 430 23071
rect 245 22999 320 23033
rect 354 22999 430 23033
rect 245 22961 430 22999
rect 245 22927 320 22961
rect 354 22927 430 22961
rect 245 22889 430 22927
rect 245 22855 320 22889
rect 354 22855 430 22889
rect 245 22817 430 22855
rect 245 22783 320 22817
rect 354 22783 430 22817
rect 245 22745 430 22783
rect 245 22711 320 22745
rect 354 22711 430 22745
rect 245 22673 430 22711
rect 245 22639 320 22673
rect 354 22639 430 22673
rect 245 22601 430 22639
rect 245 22567 320 22601
rect 354 22567 430 22601
rect 245 22529 430 22567
rect 245 22495 320 22529
rect 354 22495 430 22529
rect 245 22457 430 22495
rect 245 22423 320 22457
rect 354 22423 430 22457
rect 245 22385 430 22423
rect 245 22351 320 22385
rect 354 22351 430 22385
rect 245 22313 430 22351
rect 245 22279 320 22313
rect 354 22279 430 22313
rect 245 22241 430 22279
rect 245 22207 320 22241
rect 354 22207 430 22241
rect 245 22169 430 22207
rect 245 22135 320 22169
rect 354 22135 430 22169
rect 245 22097 430 22135
rect 245 22063 320 22097
rect 354 22063 430 22097
rect 245 22025 430 22063
rect 245 21991 320 22025
rect 354 21991 430 22025
rect 245 21953 430 21991
rect 245 21919 320 21953
rect 354 21919 430 21953
rect 245 21881 430 21919
rect 245 21847 320 21881
rect 354 21847 430 21881
rect 245 21809 430 21847
rect 245 21775 320 21809
rect 354 21775 430 21809
rect 245 21737 430 21775
rect 245 21703 320 21737
rect 354 21703 430 21737
rect 245 21665 430 21703
rect 245 21631 320 21665
rect 354 21631 430 21665
rect 245 21593 430 21631
rect 245 21559 320 21593
rect 354 21559 430 21593
rect 245 21521 430 21559
rect 245 21487 320 21521
rect 354 21487 430 21521
rect 245 21449 430 21487
rect 245 21415 320 21449
rect 354 21415 430 21449
rect 245 21377 430 21415
rect 245 21343 320 21377
rect 354 21343 430 21377
rect 245 21305 430 21343
rect 245 21271 320 21305
rect 354 21271 430 21305
rect 245 21233 430 21271
rect 245 21199 320 21233
rect 354 21199 430 21233
rect 245 21161 430 21199
rect 245 21127 320 21161
rect 354 21127 430 21161
rect 245 21089 430 21127
rect 245 21055 320 21089
rect 354 21055 430 21089
rect 245 21017 430 21055
rect 245 20983 320 21017
rect 354 20983 430 21017
rect 245 20945 430 20983
rect 245 20911 320 20945
rect 354 20911 430 20945
rect 245 20873 430 20911
rect 245 20839 320 20873
rect 354 20839 430 20873
rect 245 20801 430 20839
rect 245 20767 320 20801
rect 354 20767 430 20801
rect 245 20729 430 20767
rect 245 20695 320 20729
rect 354 20695 430 20729
rect 245 20657 430 20695
rect 245 20623 320 20657
rect 354 20623 430 20657
rect 245 20585 430 20623
rect 245 20551 320 20585
rect 354 20551 430 20585
rect 245 20513 430 20551
rect 245 20479 320 20513
rect 354 20479 430 20513
rect 245 20441 430 20479
rect 245 20407 320 20441
rect 354 20407 430 20441
rect 245 20369 430 20407
rect 245 20335 320 20369
rect 354 20335 430 20369
rect 245 20297 430 20335
rect 245 20263 320 20297
rect 354 20263 430 20297
rect 245 20225 430 20263
rect 245 20191 320 20225
rect 354 20191 430 20225
rect 245 20153 430 20191
rect 245 20119 320 20153
rect 354 20119 430 20153
rect 245 20081 430 20119
rect 245 20047 320 20081
rect 354 20047 430 20081
rect 245 20009 430 20047
rect 245 19975 320 20009
rect 354 19975 430 20009
rect 245 19937 430 19975
rect 245 19903 320 19937
rect 354 19903 430 19937
rect 245 19865 430 19903
rect 245 19831 320 19865
rect 354 19831 430 19865
rect 245 19793 430 19831
rect 245 19759 320 19793
rect 354 19759 430 19793
rect 245 19721 430 19759
rect 245 19687 320 19721
rect 354 19687 430 19721
rect 245 19649 430 19687
rect 245 19615 320 19649
rect 354 19615 430 19649
rect 245 19577 430 19615
rect 245 19543 320 19577
rect 354 19543 430 19577
rect 245 19505 430 19543
rect 245 19471 320 19505
rect 354 19471 430 19505
rect 245 19433 430 19471
rect 245 19399 320 19433
rect 354 19399 430 19433
rect 245 19361 430 19399
rect 245 19327 320 19361
rect 354 19327 430 19361
rect 245 19289 430 19327
rect 245 19255 320 19289
rect 354 19255 430 19289
rect 245 19217 430 19255
rect 245 19183 320 19217
rect 354 19183 430 19217
rect 245 19145 430 19183
rect 245 19111 320 19145
rect 354 19111 430 19145
rect 245 19073 430 19111
rect 245 19039 320 19073
rect 354 19039 430 19073
rect 245 19001 430 19039
rect 245 18967 320 19001
rect 354 18967 430 19001
rect 245 18929 430 18967
rect 245 18895 320 18929
rect 354 18895 430 18929
rect 245 18857 430 18895
rect 245 18823 320 18857
rect 354 18823 430 18857
rect 245 18785 430 18823
rect 245 18751 320 18785
rect 354 18751 430 18785
rect 245 18713 430 18751
rect 245 18679 320 18713
rect 354 18679 430 18713
rect 245 18641 430 18679
rect 245 18607 320 18641
rect 354 18607 430 18641
rect 245 18569 430 18607
rect 245 18535 320 18569
rect 354 18535 430 18569
rect 245 18497 430 18535
rect 245 18463 320 18497
rect 354 18463 430 18497
rect 245 18425 430 18463
rect 245 18391 320 18425
rect 354 18391 430 18425
rect 245 18353 430 18391
rect 245 18319 320 18353
rect 354 18319 430 18353
rect 245 18281 430 18319
rect 245 18247 320 18281
rect 354 18247 430 18281
rect 245 18209 430 18247
rect 245 18175 320 18209
rect 354 18175 430 18209
rect 245 18137 430 18175
rect 245 18103 320 18137
rect 354 18103 430 18137
rect 245 18065 430 18103
rect 245 18031 320 18065
rect 354 18031 430 18065
rect 245 17993 430 18031
rect 245 17959 320 17993
rect 354 17959 430 17993
rect 245 17921 430 17959
rect 245 17887 320 17921
rect 354 17887 430 17921
rect 245 17849 430 17887
rect 245 17815 320 17849
rect 354 17815 430 17849
rect 245 17777 430 17815
rect 245 17743 320 17777
rect 354 17743 430 17777
rect 245 17705 430 17743
rect 245 17671 320 17705
rect 354 17671 430 17705
rect 245 17633 430 17671
rect 245 17599 320 17633
rect 354 17599 430 17633
rect 245 17561 430 17599
rect 245 17527 320 17561
rect 354 17527 430 17561
rect 245 17489 430 17527
rect 245 17455 320 17489
rect 354 17455 430 17489
rect 245 17417 430 17455
rect 245 17383 320 17417
rect 354 17383 430 17417
rect 245 17345 430 17383
rect 245 17311 320 17345
rect 354 17311 430 17345
rect 245 17273 430 17311
rect 245 17239 320 17273
rect 354 17239 430 17273
rect 245 17201 430 17239
rect 245 17167 320 17201
rect 354 17167 430 17201
rect 245 17129 430 17167
rect 245 17095 320 17129
rect 354 17095 430 17129
rect 245 17057 430 17095
rect 245 17023 320 17057
rect 354 17023 430 17057
rect 245 16985 430 17023
rect 245 16951 320 16985
rect 354 16951 430 16985
rect 245 16913 430 16951
rect 245 16879 320 16913
rect 354 16879 430 16913
rect 245 16841 430 16879
rect 245 16807 320 16841
rect 354 16807 430 16841
rect 245 16769 430 16807
rect 245 16735 320 16769
rect 354 16735 430 16769
rect 245 16697 430 16735
rect 245 16663 320 16697
rect 354 16663 430 16697
rect 245 16625 430 16663
rect 245 16591 320 16625
rect 354 16591 430 16625
rect 245 16553 430 16591
rect 245 16519 320 16553
rect 354 16519 430 16553
rect 245 16481 430 16519
rect 245 16447 320 16481
rect 354 16447 430 16481
rect 245 16409 430 16447
rect 245 16375 320 16409
rect 354 16375 430 16409
rect 245 16337 430 16375
rect 245 16303 320 16337
rect 354 16303 430 16337
rect 245 16265 430 16303
rect 245 16231 320 16265
rect 354 16231 430 16265
rect 245 16193 430 16231
rect 245 16159 320 16193
rect 354 16159 430 16193
rect 245 16121 430 16159
rect 245 16087 320 16121
rect 354 16087 430 16121
rect 245 16049 430 16087
rect 245 16015 320 16049
rect 354 16015 430 16049
rect 245 15977 430 16015
rect 245 15943 320 15977
rect 354 15943 430 15977
rect 245 15905 430 15943
rect 245 15871 320 15905
rect 354 15871 430 15905
rect 245 15833 430 15871
rect 245 15799 320 15833
rect 354 15799 430 15833
rect 245 15761 430 15799
rect 245 15727 320 15761
rect 354 15727 430 15761
rect 245 15689 430 15727
rect 245 15655 320 15689
rect 354 15655 430 15689
rect 245 15617 430 15655
rect 245 15583 320 15617
rect 354 15583 430 15617
rect 245 15545 430 15583
rect 245 15511 320 15545
rect 354 15511 430 15545
rect 245 15473 430 15511
rect 245 15439 320 15473
rect 354 15439 430 15473
rect 245 15401 430 15439
rect 245 15367 320 15401
rect 354 15367 430 15401
rect 245 15329 430 15367
rect 245 15295 320 15329
rect 354 15295 430 15329
rect 245 15257 430 15295
rect 245 15223 320 15257
rect 354 15223 430 15257
rect 245 15185 430 15223
rect 245 15151 320 15185
rect 354 15151 430 15185
rect 245 15113 430 15151
rect 245 15079 320 15113
rect 354 15079 430 15113
rect 245 15041 430 15079
rect 245 15007 320 15041
rect 354 15007 430 15041
rect 245 14969 430 15007
rect 245 14935 320 14969
rect 354 14935 430 14969
tri 757 35953 760 35956 se
rect 760 35953 14216 35956
tri 14216 35953 14219 35956 sw
rect 757 35933 14219 35953
rect 757 35918 902 35933
tri 902 35918 917 35933 nw
tri 14059 35918 14074 35933 ne
rect 14074 35918 14219 35933
rect 757 35900 877 35918
rect 757 35866 807 35900
rect 841 35866 877 35900
tri 877 35893 902 35918 nw
tri 14074 35893 14099 35918 ne
rect 757 35828 877 35866
rect 757 35794 807 35828
rect 841 35794 877 35828
rect 757 35756 877 35794
rect 757 35722 807 35756
rect 841 35722 877 35756
rect 757 35684 877 35722
rect 757 35650 807 35684
rect 841 35650 877 35684
rect 757 35612 877 35650
rect 757 35578 807 35612
rect 841 35578 877 35612
rect 757 35540 877 35578
rect 757 35506 807 35540
rect 841 35506 877 35540
rect 757 35468 877 35506
rect 757 35434 807 35468
rect 841 35434 877 35468
rect 757 35396 877 35434
rect 757 35362 807 35396
rect 841 35362 877 35396
rect 757 35324 877 35362
rect 757 35290 807 35324
rect 841 35290 877 35324
rect 757 35252 877 35290
rect 757 35218 807 35252
rect 841 35218 877 35252
rect 757 35180 877 35218
rect 757 35146 807 35180
rect 841 35146 877 35180
rect 757 35108 877 35146
rect 757 35074 807 35108
rect 841 35074 877 35108
rect 757 35036 877 35074
rect 757 35002 807 35036
rect 841 35002 877 35036
rect 757 34964 877 35002
rect 757 34930 807 34964
rect 841 34930 877 34964
rect 757 34892 877 34930
rect 757 34858 807 34892
rect 841 34858 877 34892
rect 757 34820 877 34858
rect 757 34786 807 34820
rect 841 34786 877 34820
rect 757 34748 877 34786
rect 757 34714 807 34748
rect 841 34714 877 34748
rect 14099 35821 14219 35918
rect 14099 35787 14122 35821
rect 14156 35787 14219 35821
rect 14099 35749 14219 35787
rect 14099 35715 14122 35749
rect 14156 35715 14219 35749
rect 14099 35677 14219 35715
rect 14099 35643 14122 35677
rect 14156 35643 14219 35677
rect 14099 35605 14219 35643
rect 14099 35571 14122 35605
rect 14156 35571 14219 35605
rect 14099 35533 14219 35571
rect 14099 35499 14122 35533
rect 14156 35499 14219 35533
rect 14099 35461 14219 35499
rect 14099 35427 14122 35461
rect 14156 35427 14219 35461
rect 14099 35389 14219 35427
rect 14099 35355 14122 35389
rect 14156 35355 14219 35389
rect 14099 35317 14219 35355
rect 14099 35283 14122 35317
rect 14156 35283 14219 35317
rect 14099 35245 14219 35283
rect 14099 35211 14122 35245
rect 14156 35211 14219 35245
rect 14099 35173 14219 35211
rect 14099 35139 14122 35173
rect 14156 35139 14219 35173
rect 14099 35101 14219 35139
rect 14099 35067 14122 35101
rect 14156 35067 14219 35101
rect 14099 35029 14219 35067
rect 14099 34995 14122 35029
rect 14156 34995 14219 35029
rect 14099 34957 14219 34995
rect 14099 34923 14122 34957
rect 14156 34923 14219 34957
rect 14099 34885 14219 34923
rect 14099 34851 14122 34885
rect 14156 34851 14219 34885
rect 14099 34813 14219 34851
rect 14099 34779 14122 34813
rect 14156 34779 14219 34813
rect 14099 34741 14219 34779
rect 757 34676 877 34714
rect 757 34642 807 34676
rect 841 34642 877 34676
rect 757 34604 877 34642
rect 757 34570 807 34604
rect 841 34570 877 34604
rect 757 34532 877 34570
rect 757 34498 807 34532
rect 841 34498 877 34532
rect 757 34460 877 34498
rect 757 34426 807 34460
rect 841 34426 877 34460
rect 757 34388 877 34426
rect 757 34354 807 34388
rect 841 34354 877 34388
rect 757 34316 877 34354
rect 757 34282 807 34316
rect 841 34282 877 34316
rect 757 34244 877 34282
rect 757 34210 807 34244
rect 841 34210 877 34244
rect 757 34172 877 34210
rect 757 34138 807 34172
rect 841 34138 877 34172
rect 757 34100 877 34138
rect 757 34066 807 34100
rect 841 34066 877 34100
rect 757 34028 877 34066
rect 757 33994 807 34028
rect 841 33994 877 34028
rect 757 33956 877 33994
rect 757 33922 807 33956
rect 841 33922 877 33956
rect 757 33884 877 33922
rect 757 33850 807 33884
rect 841 33850 877 33884
rect 757 33812 877 33850
rect 757 33778 807 33812
rect 841 33778 877 33812
rect 757 33740 877 33778
rect 757 33706 807 33740
rect 841 33706 877 33740
rect 757 33668 877 33706
rect 757 33634 807 33668
rect 841 33634 877 33668
rect 757 33596 877 33634
rect 757 33562 807 33596
rect 841 33562 877 33596
rect 757 33524 877 33562
rect 757 33490 807 33524
rect 841 33490 877 33524
rect 757 33452 877 33490
rect 757 33418 807 33452
rect 841 33418 877 33452
rect 757 33380 877 33418
rect 757 33346 807 33380
rect 841 33346 877 33380
rect 757 33308 877 33346
rect 757 33274 807 33308
rect 841 33274 877 33308
rect 757 33236 877 33274
rect 757 33202 807 33236
rect 841 33202 877 33236
rect 757 33164 877 33202
rect 757 33130 807 33164
rect 841 33130 877 33164
rect 757 33092 877 33130
rect 757 33058 807 33092
rect 841 33058 877 33092
rect 757 33020 877 33058
rect 757 32986 807 33020
rect 841 32986 877 33020
rect 757 32948 877 32986
rect 757 32914 807 32948
rect 841 32914 877 32948
rect 757 32876 877 32914
rect 757 32842 807 32876
rect 841 32842 877 32876
rect 757 32804 877 32842
rect 757 32770 807 32804
rect 841 32770 877 32804
rect 757 32732 877 32770
rect 757 32698 807 32732
rect 841 32698 877 32732
rect 757 32660 877 32698
rect 757 32626 807 32660
rect 841 32626 877 32660
rect 757 32588 877 32626
rect 757 32554 807 32588
rect 841 32554 877 32588
rect 757 32516 877 32554
rect 757 32482 807 32516
rect 841 32482 877 32516
rect 757 32444 877 32482
rect 757 32410 807 32444
rect 841 32410 877 32444
rect 757 32372 877 32410
rect 757 32338 807 32372
rect 841 32338 877 32372
rect 757 32300 877 32338
rect 757 32266 807 32300
rect 841 32266 877 32300
rect 757 32228 877 32266
rect 757 32194 807 32228
rect 841 32194 877 32228
rect 757 32156 877 32194
rect 757 32122 807 32156
rect 841 32122 877 32156
rect 757 32084 877 32122
rect 757 32050 807 32084
rect 841 32050 877 32084
rect 757 32012 877 32050
rect 757 31978 807 32012
rect 841 31978 877 32012
rect 757 31940 877 31978
rect 757 31906 807 31940
rect 841 31906 877 31940
rect 757 31868 877 31906
rect 757 31834 807 31868
rect 841 31834 877 31868
rect 757 31796 877 31834
rect 757 31762 807 31796
rect 841 31762 877 31796
rect 757 31724 877 31762
rect 757 31690 807 31724
rect 841 31690 877 31724
rect 757 31652 877 31690
rect 757 31618 807 31652
rect 841 31618 877 31652
rect 757 31580 877 31618
rect 757 31546 807 31580
rect 841 31546 877 31580
rect 757 31508 877 31546
rect 757 31474 807 31508
rect 841 31474 877 31508
rect 757 31436 877 31474
rect 757 31402 807 31436
rect 841 31402 877 31436
rect 757 31364 877 31402
rect 757 31330 807 31364
rect 841 31330 877 31364
rect 757 31292 877 31330
rect 757 31258 807 31292
rect 841 31258 877 31292
rect 757 31220 877 31258
rect 757 31186 807 31220
rect 841 31186 877 31220
rect 757 31148 877 31186
rect 757 31114 807 31148
rect 841 31114 877 31148
rect 757 31076 877 31114
rect 757 31042 807 31076
rect 841 31042 877 31076
rect 757 31004 877 31042
rect 757 30970 807 31004
rect 841 30970 877 31004
rect 757 30932 877 30970
rect 757 30898 807 30932
rect 841 30898 877 30932
rect 757 30860 877 30898
rect 757 30826 807 30860
rect 841 30826 877 30860
rect 757 30788 877 30826
rect 757 30754 807 30788
rect 841 30754 877 30788
rect 757 30716 877 30754
rect 757 30682 807 30716
rect 841 30682 877 30716
rect 757 30644 877 30682
rect 757 30610 807 30644
rect 841 30610 877 30644
rect 757 30572 877 30610
rect 757 30538 807 30572
rect 841 30538 877 30572
rect 757 30500 877 30538
rect 757 30466 807 30500
rect 841 30466 877 30500
rect 757 30428 877 30466
rect 757 30394 807 30428
rect 841 30394 877 30428
rect 757 30356 877 30394
rect 757 30322 807 30356
rect 841 30322 877 30356
rect 757 30284 877 30322
rect 757 30250 807 30284
rect 841 30250 877 30284
rect 757 30212 877 30250
rect 757 30178 807 30212
rect 841 30178 877 30212
rect 757 30140 877 30178
rect 757 30106 807 30140
rect 841 30106 877 30140
rect 757 30068 877 30106
rect 757 30034 807 30068
rect 841 30034 877 30068
rect 757 29996 877 30034
rect 757 29962 807 29996
rect 841 29962 877 29996
rect 757 29924 877 29962
rect 757 29890 807 29924
rect 841 29890 877 29924
rect 757 29852 877 29890
rect 757 29818 807 29852
rect 841 29818 877 29852
rect 757 29780 877 29818
rect 757 29746 807 29780
rect 841 29746 877 29780
rect 757 29708 877 29746
rect 757 29674 807 29708
rect 841 29674 877 29708
rect 757 29636 877 29674
rect 757 29602 807 29636
rect 841 29602 877 29636
rect 757 29564 877 29602
rect 757 29530 807 29564
rect 841 29530 877 29564
rect 757 29492 877 29530
rect 757 29458 807 29492
rect 841 29458 877 29492
rect 757 29420 877 29458
rect 757 29386 807 29420
rect 841 29386 877 29420
rect 757 29348 877 29386
rect 757 29314 807 29348
rect 841 29314 877 29348
rect 757 29276 877 29314
rect 757 29242 807 29276
rect 841 29242 877 29276
rect 757 29204 877 29242
rect 757 29170 807 29204
rect 841 29170 877 29204
rect 757 29132 877 29170
rect 757 29098 807 29132
rect 841 29098 877 29132
rect 757 29060 877 29098
rect 757 29026 807 29060
rect 841 29026 877 29060
rect 757 28988 877 29026
rect 757 28954 807 28988
rect 841 28954 877 28988
rect 757 28916 877 28954
rect 757 28882 807 28916
rect 841 28882 877 28916
rect 757 28844 877 28882
rect 757 28810 807 28844
rect 841 28810 877 28844
rect 757 28772 877 28810
rect 757 28738 807 28772
rect 841 28738 877 28772
rect 757 28700 877 28738
rect 757 28666 807 28700
rect 841 28666 877 28700
rect 757 28628 877 28666
rect 757 28594 807 28628
rect 841 28594 877 28628
rect 757 28556 877 28594
rect 757 28522 807 28556
rect 841 28522 877 28556
rect 757 28484 877 28522
rect 757 28450 807 28484
rect 841 28450 877 28484
rect 757 28412 877 28450
rect 757 28378 807 28412
rect 841 28378 877 28412
rect 757 28340 877 28378
rect 757 28306 807 28340
rect 841 28306 877 28340
rect 757 28268 877 28306
rect 757 28234 807 28268
rect 841 28234 877 28268
rect 757 28196 877 28234
rect 757 28162 807 28196
rect 841 28162 877 28196
rect 757 28124 877 28162
rect 757 28090 807 28124
rect 841 28090 877 28124
rect 757 28052 877 28090
rect 757 28018 807 28052
rect 841 28018 877 28052
rect 757 27980 877 28018
rect 757 27946 807 27980
rect 841 27946 877 27980
rect 757 27908 877 27946
rect 757 27874 807 27908
rect 841 27874 877 27908
rect 757 27836 877 27874
rect 757 27802 807 27836
rect 841 27802 877 27836
rect 757 27764 877 27802
rect 757 27730 807 27764
rect 841 27730 877 27764
rect 757 27692 877 27730
rect 757 27658 807 27692
rect 841 27658 877 27692
rect 757 27620 877 27658
rect 757 27586 807 27620
rect 841 27586 877 27620
rect 757 27548 877 27586
rect 757 27514 807 27548
rect 841 27514 877 27548
rect 757 27476 877 27514
rect 757 27442 807 27476
rect 841 27442 877 27476
rect 757 27404 877 27442
rect 757 27370 807 27404
rect 841 27370 877 27404
rect 757 27332 877 27370
rect 757 27298 807 27332
rect 841 27298 877 27332
rect 757 27260 877 27298
rect 757 27226 807 27260
rect 841 27226 877 27260
rect 757 27188 877 27226
rect 757 27154 807 27188
rect 841 27154 877 27188
rect 757 27116 877 27154
rect 757 27082 807 27116
rect 841 27082 877 27116
rect 757 27044 877 27082
rect 757 27010 807 27044
rect 841 27010 877 27044
rect 757 26972 877 27010
rect 757 26938 807 26972
rect 841 26938 877 26972
rect 757 26900 877 26938
rect 757 26866 807 26900
rect 841 26866 877 26900
rect 757 26828 877 26866
rect 757 26794 807 26828
rect 841 26794 877 26828
rect 757 26756 877 26794
rect 757 26722 807 26756
rect 841 26722 877 26756
rect 757 26684 877 26722
rect 757 26650 807 26684
rect 841 26650 877 26684
rect 757 26612 877 26650
rect 757 26578 807 26612
rect 841 26578 877 26612
rect 757 26540 877 26578
rect 757 26506 807 26540
rect 841 26506 877 26540
rect 757 26468 877 26506
rect 757 26434 807 26468
rect 841 26434 877 26468
rect 757 26396 877 26434
rect 757 26362 807 26396
rect 841 26362 877 26396
rect 757 26324 877 26362
rect 757 26290 807 26324
rect 841 26290 877 26324
rect 757 26252 877 26290
rect 757 26218 807 26252
rect 841 26218 877 26252
rect 757 26180 877 26218
rect 757 26146 807 26180
rect 841 26146 877 26180
rect 757 26108 877 26146
rect 757 26074 807 26108
rect 841 26074 877 26108
rect 757 26036 877 26074
rect 757 26002 807 26036
rect 841 26002 877 26036
rect 757 25964 877 26002
rect 757 25930 807 25964
rect 841 25930 877 25964
rect 757 25892 877 25930
rect 757 25858 807 25892
rect 841 25858 877 25892
rect 757 25820 877 25858
rect 757 25786 807 25820
rect 841 25786 877 25820
rect 757 25748 877 25786
rect 757 25714 807 25748
rect 841 25714 877 25748
rect 757 25676 877 25714
rect 757 25642 807 25676
rect 841 25642 877 25676
rect 757 25604 877 25642
rect 757 25570 807 25604
rect 841 25570 877 25604
rect 757 25532 877 25570
rect 757 25498 807 25532
rect 841 25498 877 25532
rect 757 25460 877 25498
rect 757 25426 807 25460
rect 841 25426 877 25460
rect 757 25388 877 25426
rect 757 25354 807 25388
rect 841 25354 877 25388
rect 757 25316 877 25354
rect 757 25282 807 25316
rect 841 25282 877 25316
rect 757 25244 877 25282
rect 757 25210 807 25244
rect 841 25210 877 25244
rect 757 25172 877 25210
rect 757 25138 807 25172
rect 841 25138 877 25172
rect 757 25100 877 25138
rect 757 25066 807 25100
rect 841 25066 877 25100
rect 757 25028 877 25066
rect 757 24994 807 25028
rect 841 24994 877 25028
rect 757 24956 877 24994
rect 757 24922 807 24956
rect 841 24922 877 24956
rect 757 24884 877 24922
rect 757 24850 807 24884
rect 841 24850 877 24884
rect 757 24812 877 24850
rect 757 24778 807 24812
rect 841 24778 877 24812
rect 757 24740 877 24778
rect 757 24706 807 24740
rect 841 24706 877 24740
rect 757 24668 877 24706
rect 757 24634 807 24668
rect 841 24634 877 24668
rect 757 24596 877 24634
rect 757 24562 807 24596
rect 841 24562 877 24596
rect 757 24524 877 24562
rect 757 24490 807 24524
rect 841 24490 877 24524
rect 757 24452 877 24490
rect 757 24418 807 24452
rect 841 24418 877 24452
rect 757 24380 877 24418
rect 757 24346 807 24380
rect 841 24346 877 24380
rect 757 24308 877 24346
rect 757 24274 807 24308
rect 841 24274 877 24308
rect 757 24236 877 24274
rect 757 24202 807 24236
rect 841 24202 877 24236
rect 757 24164 877 24202
rect 757 24130 807 24164
rect 841 24130 877 24164
rect 757 24092 877 24130
rect 757 24058 807 24092
rect 841 24058 877 24092
rect 757 24020 877 24058
rect 757 23986 807 24020
rect 841 23986 877 24020
rect 757 23948 877 23986
rect 757 23914 807 23948
rect 841 23914 877 23948
rect 757 23876 877 23914
rect 757 23842 807 23876
rect 841 23842 877 23876
rect 757 23804 877 23842
rect 757 23770 807 23804
rect 841 23770 877 23804
rect 757 23732 877 23770
rect 757 23698 807 23732
rect 841 23698 877 23732
rect 757 23660 877 23698
rect 757 23626 807 23660
rect 841 23626 877 23660
rect 757 23588 877 23626
rect 757 23554 807 23588
rect 841 23554 877 23588
rect 757 23516 877 23554
rect 757 23482 807 23516
rect 841 23482 877 23516
rect 757 23444 877 23482
rect 757 23410 807 23444
rect 841 23410 877 23444
rect 757 23372 877 23410
rect 757 23338 807 23372
rect 841 23338 877 23372
rect 757 23300 877 23338
rect 757 23266 807 23300
rect 841 23266 877 23300
rect 757 23228 877 23266
rect 757 23194 807 23228
rect 841 23194 877 23228
rect 757 23156 877 23194
rect 757 23122 807 23156
rect 841 23122 877 23156
rect 757 23084 877 23122
rect 757 23050 807 23084
rect 841 23050 877 23084
rect 757 23012 877 23050
rect 757 22978 807 23012
rect 841 22978 877 23012
rect 757 22940 877 22978
rect 757 22906 807 22940
rect 841 22906 877 22940
rect 757 22868 877 22906
rect 757 22834 807 22868
rect 841 22834 877 22868
rect 757 22796 877 22834
rect 757 22762 807 22796
rect 841 22762 877 22796
rect 757 22724 877 22762
rect 757 22690 807 22724
rect 841 22690 877 22724
rect 757 22652 877 22690
rect 757 22618 807 22652
rect 841 22618 877 22652
rect 757 22580 877 22618
rect 757 22546 807 22580
rect 841 22546 877 22580
rect 757 22508 877 22546
rect 757 22474 807 22508
rect 841 22474 877 22508
rect 757 22436 877 22474
rect 757 22402 807 22436
rect 841 22402 877 22436
rect 757 22364 877 22402
rect 757 22330 807 22364
rect 841 22330 877 22364
rect 757 22292 877 22330
rect 757 22258 807 22292
rect 841 22258 877 22292
rect 757 22220 877 22258
rect 757 22186 807 22220
rect 841 22186 877 22220
rect 757 22148 877 22186
rect 757 22114 807 22148
rect 841 22114 877 22148
rect 757 22076 877 22114
rect 757 22042 807 22076
rect 841 22042 877 22076
rect 757 22004 877 22042
rect 757 21970 807 22004
rect 841 21970 877 22004
rect 757 21932 877 21970
rect 757 21898 807 21932
rect 841 21898 877 21932
rect 757 21860 877 21898
rect 757 21826 807 21860
rect 841 21826 877 21860
rect 757 21788 877 21826
rect 757 21754 807 21788
rect 841 21754 877 21788
rect 757 21716 877 21754
rect 757 21682 807 21716
rect 841 21682 877 21716
rect 757 21644 877 21682
rect 757 21610 807 21644
rect 841 21610 877 21644
rect 757 21572 877 21610
rect 757 21538 807 21572
rect 841 21538 877 21572
rect 757 21500 877 21538
rect 757 21466 807 21500
rect 841 21466 877 21500
rect 757 21428 877 21466
rect 757 21394 807 21428
rect 841 21394 877 21428
rect 757 21356 877 21394
rect 757 21322 807 21356
rect 841 21322 877 21356
rect 757 21284 877 21322
rect 757 21250 807 21284
rect 841 21250 877 21284
rect 757 21212 877 21250
rect 757 21178 807 21212
rect 841 21178 877 21212
rect 757 21140 877 21178
rect 757 21106 807 21140
rect 841 21106 877 21140
rect 757 21068 877 21106
rect 757 21034 807 21068
rect 841 21034 877 21068
rect 757 20996 877 21034
rect 757 20962 807 20996
rect 841 20962 877 20996
rect 757 20924 877 20962
rect 757 20890 807 20924
rect 841 20890 877 20924
rect 757 20852 877 20890
rect 757 20818 807 20852
rect 841 20818 877 20852
rect 757 20780 877 20818
rect 757 20746 807 20780
rect 841 20746 877 20780
rect 757 20708 877 20746
rect 757 20674 807 20708
rect 841 20674 877 20708
rect 757 20636 877 20674
rect 757 20602 807 20636
rect 841 20602 877 20636
rect 757 20564 877 20602
rect 757 20530 807 20564
rect 841 20530 877 20564
rect 757 20492 877 20530
rect 757 20458 807 20492
rect 841 20458 877 20492
rect 757 20420 877 20458
rect 757 20386 807 20420
rect 841 20386 877 20420
rect 757 20348 877 20386
rect 757 20314 807 20348
rect 841 20314 877 20348
rect 757 20276 877 20314
rect 757 20242 807 20276
rect 841 20242 877 20276
rect 757 20204 877 20242
rect 757 20170 807 20204
rect 841 20170 877 20204
rect 757 20132 877 20170
rect 757 20098 807 20132
rect 841 20098 877 20132
rect 757 20060 877 20098
rect 757 20026 807 20060
rect 841 20026 877 20060
rect 757 19988 877 20026
rect 757 19954 807 19988
rect 841 19954 877 19988
rect 757 19916 877 19954
rect 757 19882 807 19916
rect 841 19882 877 19916
rect 757 19844 877 19882
rect 757 19810 807 19844
rect 841 19810 877 19844
rect 757 19772 877 19810
rect 757 19738 807 19772
rect 841 19738 877 19772
rect 757 19700 877 19738
rect 757 19666 807 19700
rect 841 19666 877 19700
rect 757 19628 877 19666
rect 757 19594 807 19628
rect 841 19594 877 19628
rect 757 19556 877 19594
rect 757 19522 807 19556
rect 841 19522 877 19556
rect 757 19484 877 19522
rect 757 19450 807 19484
rect 841 19450 877 19484
rect 757 19412 877 19450
rect 757 19378 807 19412
rect 841 19378 877 19412
rect 757 19340 877 19378
rect 757 19306 807 19340
rect 841 19306 877 19340
rect 757 19268 877 19306
rect 757 19234 807 19268
rect 841 19234 877 19268
rect 757 19196 877 19234
rect 757 19162 807 19196
rect 841 19162 877 19196
rect 757 19124 877 19162
rect 757 19090 807 19124
rect 841 19090 877 19124
rect 757 19052 877 19090
rect 757 19018 807 19052
rect 841 19018 877 19052
rect 757 18980 877 19018
rect 757 18946 807 18980
rect 841 18946 877 18980
rect 757 18908 877 18946
rect 757 18874 807 18908
rect 841 18874 877 18908
rect 757 18836 877 18874
rect 757 18802 807 18836
rect 841 18802 877 18836
rect 757 18764 877 18802
rect 757 18730 807 18764
rect 841 18730 877 18764
rect 757 18692 877 18730
rect 757 18658 807 18692
rect 841 18658 877 18692
rect 757 18620 877 18658
rect 757 18586 807 18620
rect 841 18586 877 18620
rect 757 18548 877 18586
rect 757 18514 807 18548
rect 841 18514 877 18548
rect 757 18476 877 18514
rect 757 18442 807 18476
rect 841 18442 877 18476
rect 757 18404 877 18442
rect 757 18370 807 18404
rect 841 18370 877 18404
rect 757 18332 877 18370
rect 757 18298 807 18332
rect 841 18298 877 18332
rect 757 18260 877 18298
rect 757 18226 807 18260
rect 841 18226 877 18260
rect 757 18188 877 18226
rect 757 18154 807 18188
rect 841 18154 877 18188
rect 757 18116 877 18154
rect 757 18082 807 18116
rect 841 18082 877 18116
rect 757 18044 877 18082
rect 757 18010 807 18044
rect 841 18010 877 18044
rect 757 17972 877 18010
rect 757 17938 807 17972
rect 841 17938 877 17972
rect 757 17900 877 17938
rect 757 17866 807 17900
rect 841 17866 877 17900
rect 757 17828 877 17866
rect 757 17794 807 17828
rect 841 17794 877 17828
rect 757 17756 877 17794
rect 757 17722 807 17756
rect 841 17722 877 17756
rect 757 17684 877 17722
rect 757 17650 807 17684
rect 841 17650 877 17684
rect 757 17612 877 17650
rect 757 17578 807 17612
rect 841 17578 877 17612
rect 757 17540 877 17578
rect 757 17506 807 17540
rect 841 17506 877 17540
rect 757 17468 877 17506
rect 757 17434 807 17468
rect 841 17434 877 17468
rect 757 17396 877 17434
rect 757 17362 807 17396
rect 841 17362 877 17396
rect 757 17324 877 17362
rect 757 17290 807 17324
rect 841 17290 877 17324
rect 757 17252 877 17290
rect 757 17218 807 17252
rect 841 17218 877 17252
rect 757 17180 877 17218
rect 757 17146 807 17180
rect 841 17146 877 17180
rect 757 17108 877 17146
rect 757 17074 807 17108
rect 841 17074 877 17108
rect 757 17036 877 17074
rect 757 17002 807 17036
rect 841 17002 877 17036
rect 757 16964 877 17002
rect 757 16930 807 16964
rect 841 16930 877 16964
rect 757 16892 877 16930
rect 757 16858 807 16892
rect 841 16858 877 16892
rect 757 16820 877 16858
rect 757 16786 807 16820
rect 841 16786 877 16820
rect 757 16748 877 16786
rect 757 16714 807 16748
rect 841 16714 877 16748
rect 757 16676 877 16714
rect 757 16642 807 16676
rect 841 16642 877 16676
rect 757 16604 877 16642
rect 757 16570 807 16604
rect 841 16570 877 16604
rect 757 16532 877 16570
rect 757 16498 807 16532
rect 841 16498 877 16532
rect 757 16460 877 16498
rect 757 16426 807 16460
rect 841 16426 877 16460
rect 757 16388 877 16426
rect 757 16354 807 16388
rect 841 16354 877 16388
rect 757 16316 877 16354
rect 757 16282 807 16316
rect 841 16282 877 16316
rect 757 16244 877 16282
rect 757 16210 807 16244
rect 841 16210 877 16244
rect 757 16172 877 16210
rect 757 16138 807 16172
rect 841 16138 877 16172
rect 757 16100 877 16138
rect 757 16066 807 16100
rect 841 16066 877 16100
rect 757 16028 877 16066
rect 757 15994 807 16028
rect 841 15994 877 16028
rect 757 15956 877 15994
rect 757 15922 807 15956
rect 841 15922 877 15956
rect 757 15884 877 15922
rect 757 15850 807 15884
rect 841 15850 877 15884
rect 757 15812 877 15850
rect 757 15778 807 15812
rect 841 15778 877 15812
rect 757 15740 877 15778
rect 757 15706 807 15740
rect 841 15706 877 15740
rect 757 15668 877 15706
rect 757 15634 807 15668
rect 841 15634 877 15668
rect 757 15596 877 15634
rect 757 15562 807 15596
rect 841 15562 877 15596
rect 757 15524 877 15562
rect 757 15490 807 15524
rect 841 15490 877 15524
rect 757 15452 877 15490
rect 757 15418 807 15452
rect 841 15418 877 15452
rect 757 15380 877 15418
rect 757 15346 807 15380
rect 841 15346 877 15380
rect 757 15308 877 15346
rect 757 15274 807 15308
rect 841 15274 877 15308
rect 757 15236 877 15274
rect 757 15202 807 15236
rect 841 15202 877 15236
rect 757 15164 877 15202
rect 1119 34679 13887 34721
rect 1119 34645 1301 34679
rect 1335 34645 1373 34679
rect 1407 34645 1445 34679
rect 1479 34645 1517 34679
rect 1551 34645 1589 34679
rect 1623 34645 1661 34679
rect 1695 34645 1733 34679
rect 1767 34645 1805 34679
rect 1839 34645 1877 34679
rect 1911 34645 1949 34679
rect 1983 34645 2021 34679
rect 2055 34645 2093 34679
rect 2127 34645 2165 34679
rect 2199 34645 2237 34679
rect 2271 34645 2309 34679
rect 2343 34645 2381 34679
rect 2415 34645 2453 34679
rect 2487 34645 2525 34679
rect 2559 34645 2597 34679
rect 2631 34645 2669 34679
rect 2703 34645 2741 34679
rect 2775 34645 2813 34679
rect 2847 34645 2885 34679
rect 2919 34645 2957 34679
rect 2991 34645 3029 34679
rect 3063 34645 3101 34679
rect 3135 34645 3173 34679
rect 3207 34645 3245 34679
rect 3279 34645 3317 34679
rect 3351 34645 3389 34679
rect 3423 34645 3461 34679
rect 3495 34645 3533 34679
rect 3567 34645 3605 34679
rect 3639 34645 3677 34679
rect 3711 34645 3749 34679
rect 3783 34645 3821 34679
rect 3855 34645 3893 34679
rect 3927 34645 3965 34679
rect 3999 34645 4037 34679
rect 4071 34645 4109 34679
rect 4143 34645 4181 34679
rect 4215 34645 4253 34679
rect 4287 34645 4325 34679
rect 4359 34645 4397 34679
rect 4431 34645 4469 34679
rect 4503 34645 4541 34679
rect 4575 34645 4613 34679
rect 4647 34645 4685 34679
rect 4719 34645 4757 34679
rect 4791 34645 4829 34679
rect 4863 34645 4901 34679
rect 4935 34645 4973 34679
rect 5007 34645 5045 34679
rect 5079 34645 5117 34679
rect 5151 34645 5189 34679
rect 5223 34645 5261 34679
rect 5295 34645 5333 34679
rect 5367 34645 5405 34679
rect 5439 34645 5477 34679
rect 5511 34645 5549 34679
rect 5583 34645 5621 34679
rect 5655 34645 5693 34679
rect 5727 34645 5765 34679
rect 5799 34645 5837 34679
rect 5871 34645 5909 34679
rect 5943 34645 5981 34679
rect 6015 34645 6053 34679
rect 6087 34645 6125 34679
rect 6159 34645 6197 34679
rect 6231 34645 6269 34679
rect 6303 34645 6341 34679
rect 6375 34645 6413 34679
rect 6447 34645 6485 34679
rect 6519 34645 6557 34679
rect 6591 34645 6629 34679
rect 6663 34645 6701 34679
rect 6735 34645 6773 34679
rect 6807 34645 6845 34679
rect 6879 34645 6917 34679
rect 6951 34645 6989 34679
rect 7023 34645 7061 34679
rect 7095 34645 7133 34679
rect 7167 34645 7205 34679
rect 7239 34645 7277 34679
rect 7311 34645 7349 34679
rect 7383 34645 7421 34679
rect 7455 34645 7493 34679
rect 7527 34645 7565 34679
rect 7599 34645 7637 34679
rect 7671 34645 7709 34679
rect 7743 34645 7781 34679
rect 7815 34645 7853 34679
rect 7887 34645 7925 34679
rect 7959 34645 7997 34679
rect 8031 34645 8069 34679
rect 8103 34645 8141 34679
rect 8175 34645 8213 34679
rect 8247 34645 8285 34679
rect 8319 34645 8357 34679
rect 8391 34645 8429 34679
rect 8463 34645 8501 34679
rect 8535 34645 8573 34679
rect 8607 34645 8645 34679
rect 8679 34645 8717 34679
rect 8751 34645 8789 34679
rect 8823 34645 8861 34679
rect 8895 34645 8933 34679
rect 8967 34645 9005 34679
rect 9039 34645 9077 34679
rect 9111 34645 9149 34679
rect 9183 34645 9221 34679
rect 9255 34645 9293 34679
rect 9327 34645 9365 34679
rect 9399 34645 9437 34679
rect 9471 34645 9509 34679
rect 9543 34645 9581 34679
rect 9615 34645 9653 34679
rect 9687 34645 9725 34679
rect 9759 34645 9797 34679
rect 9831 34645 9869 34679
rect 9903 34645 9941 34679
rect 9975 34645 10013 34679
rect 10047 34645 10085 34679
rect 10119 34645 10157 34679
rect 10191 34645 10229 34679
rect 10263 34645 10301 34679
rect 10335 34645 10373 34679
rect 10407 34645 10445 34679
rect 10479 34645 10517 34679
rect 10551 34645 10589 34679
rect 10623 34645 10661 34679
rect 10695 34645 10733 34679
rect 10767 34645 10805 34679
rect 10839 34645 10877 34679
rect 10911 34645 10949 34679
rect 10983 34645 11021 34679
rect 11055 34645 11093 34679
rect 11127 34645 11165 34679
rect 11199 34645 11237 34679
rect 11271 34645 11309 34679
rect 11343 34645 11381 34679
rect 11415 34645 11453 34679
rect 11487 34645 11525 34679
rect 11559 34645 11597 34679
rect 11631 34645 11669 34679
rect 11703 34645 11741 34679
rect 11775 34645 11813 34679
rect 11847 34645 11885 34679
rect 11919 34645 11957 34679
rect 11991 34645 12029 34679
rect 12063 34645 12101 34679
rect 12135 34645 12173 34679
rect 12207 34645 12245 34679
rect 12279 34645 12317 34679
rect 12351 34645 12389 34679
rect 12423 34645 12461 34679
rect 12495 34645 12533 34679
rect 12567 34645 12605 34679
rect 12639 34645 12677 34679
rect 12711 34645 12749 34679
rect 12783 34645 12821 34679
rect 12855 34645 12893 34679
rect 12927 34645 12965 34679
rect 12999 34645 13037 34679
rect 13071 34645 13109 34679
rect 13143 34645 13181 34679
rect 13215 34645 13253 34679
rect 13287 34645 13325 34679
rect 13359 34645 13397 34679
rect 13431 34645 13469 34679
rect 13503 34645 13541 34679
rect 13575 34645 13613 34679
rect 13647 34645 13685 34679
rect 13719 34645 13887 34679
rect 1119 34603 13887 34645
rect 1119 34482 1237 34603
rect 1119 34448 1161 34482
rect 1195 34448 1237 34482
rect 1119 34410 1237 34448
rect 1119 34376 1161 34410
rect 1195 34376 1237 34410
rect 1119 34338 1237 34376
rect 1119 34304 1161 34338
rect 1195 34304 1237 34338
rect 1119 34266 1237 34304
rect 1119 34232 1161 34266
rect 1195 34232 1237 34266
rect 1119 34194 1237 34232
rect 1119 34160 1161 34194
rect 1195 34160 1237 34194
rect 1119 34122 1237 34160
rect 1119 34088 1161 34122
rect 1195 34088 1237 34122
rect 1119 34050 1237 34088
rect 1119 34016 1161 34050
rect 1195 34016 1237 34050
rect 1119 33978 1237 34016
rect 1119 33944 1161 33978
rect 1195 33944 1237 33978
rect 1119 33906 1237 33944
rect 1119 33872 1161 33906
rect 1195 33872 1237 33906
rect 1119 33834 1237 33872
rect 1119 33800 1161 33834
rect 1195 33800 1237 33834
rect 1119 33762 1237 33800
rect 1119 33728 1161 33762
rect 1195 33728 1237 33762
rect 1119 33690 1237 33728
rect 1119 33656 1161 33690
rect 1195 33656 1237 33690
rect 1119 33618 1237 33656
rect 1119 33584 1161 33618
rect 1195 33584 1237 33618
rect 1119 33546 1237 33584
rect 1119 33512 1161 33546
rect 1195 33512 1237 33546
rect 1119 33474 1237 33512
rect 1119 33440 1161 33474
rect 1195 33440 1237 33474
rect 1119 33402 1237 33440
rect 1119 33368 1161 33402
rect 1195 33368 1237 33402
rect 1119 33330 1237 33368
rect 1119 33296 1161 33330
rect 1195 33296 1237 33330
rect 1119 33258 1237 33296
rect 1119 33224 1161 33258
rect 1195 33224 1237 33258
rect 1119 33186 1237 33224
rect 1119 33152 1161 33186
rect 1195 33152 1237 33186
rect 1119 33114 1237 33152
rect 1119 33080 1161 33114
rect 1195 33080 1237 33114
rect 1119 33042 1237 33080
rect 1119 33008 1161 33042
rect 1195 33008 1237 33042
rect 1119 32970 1237 33008
rect 1119 32936 1161 32970
rect 1195 32936 1237 32970
rect 1119 32898 1237 32936
rect 1119 32864 1161 32898
rect 1195 32864 1237 32898
rect 1119 32826 1237 32864
rect 1119 32792 1161 32826
rect 1195 32792 1237 32826
rect 1119 32754 1237 32792
rect 1119 32720 1161 32754
rect 1195 32720 1237 32754
rect 1119 32682 1237 32720
rect 1119 32648 1161 32682
rect 1195 32648 1237 32682
rect 1119 32610 1237 32648
rect 1119 32576 1161 32610
rect 1195 32576 1237 32610
rect 1119 32538 1237 32576
rect 1119 32504 1161 32538
rect 1195 32504 1237 32538
rect 1119 32466 1237 32504
rect 1119 32432 1161 32466
rect 1195 32432 1237 32466
rect 1119 32394 1237 32432
rect 1119 32360 1161 32394
rect 1195 32360 1237 32394
rect 1119 32322 1237 32360
rect 1119 32288 1161 32322
rect 1195 32288 1237 32322
rect 1119 32250 1237 32288
rect 1119 32216 1161 32250
rect 1195 32216 1237 32250
rect 1119 32178 1237 32216
rect 1119 32144 1161 32178
rect 1195 32144 1237 32178
rect 1119 32106 1237 32144
rect 1119 32072 1161 32106
rect 1195 32072 1237 32106
rect 1119 32034 1237 32072
rect 1119 32000 1161 32034
rect 1195 32000 1237 32034
rect 1119 31962 1237 32000
rect 1119 31928 1161 31962
rect 1195 31928 1237 31962
rect 1119 31890 1237 31928
rect 1119 31856 1161 31890
rect 1195 31856 1237 31890
rect 1119 31818 1237 31856
rect 1119 31784 1161 31818
rect 1195 31784 1237 31818
rect 1119 31746 1237 31784
rect 1119 31712 1161 31746
rect 1195 31712 1237 31746
rect 1119 31674 1237 31712
rect 1119 31640 1161 31674
rect 1195 31640 1237 31674
rect 1119 31602 1237 31640
rect 1119 31568 1161 31602
rect 1195 31568 1237 31602
rect 1119 31530 1237 31568
rect 1119 31496 1161 31530
rect 1195 31496 1237 31530
rect 1119 31458 1237 31496
rect 1119 31424 1161 31458
rect 1195 31424 1237 31458
rect 1119 31386 1237 31424
rect 1119 31352 1161 31386
rect 1195 31352 1237 31386
rect 1119 31314 1237 31352
rect 1119 31280 1161 31314
rect 1195 31280 1237 31314
rect 1119 31242 1237 31280
rect 1119 31208 1161 31242
rect 1195 31208 1237 31242
rect 1119 31170 1237 31208
rect 1119 31136 1161 31170
rect 1195 31136 1237 31170
rect 1119 31098 1237 31136
rect 1119 31064 1161 31098
rect 1195 31064 1237 31098
rect 1119 31026 1237 31064
rect 1119 30992 1161 31026
rect 1195 30992 1237 31026
rect 1119 30954 1237 30992
rect 1119 30920 1161 30954
rect 1195 30920 1237 30954
rect 1119 30882 1237 30920
rect 1119 30848 1161 30882
rect 1195 30848 1237 30882
rect 1119 30810 1237 30848
rect 1119 30776 1161 30810
rect 1195 30776 1237 30810
rect 1119 30738 1237 30776
rect 1119 30704 1161 30738
rect 1195 30704 1237 30738
rect 1119 30666 1237 30704
rect 1119 30632 1161 30666
rect 1195 30632 1237 30666
rect 1119 30594 1237 30632
rect 1119 30560 1161 30594
rect 1195 30560 1237 30594
rect 1119 30522 1237 30560
rect 1119 30488 1161 30522
rect 1195 30488 1237 30522
rect 1119 30450 1237 30488
rect 1119 30416 1161 30450
rect 1195 30416 1237 30450
rect 1119 30378 1237 30416
rect 1119 30344 1161 30378
rect 1195 30344 1237 30378
rect 1119 30306 1237 30344
rect 1119 30272 1161 30306
rect 1195 30281 1237 30306
rect 13769 34474 13887 34603
rect 13769 34440 13809 34474
rect 13843 34440 13887 34474
rect 13769 34402 13887 34440
rect 13769 34368 13809 34402
rect 13843 34368 13887 34402
rect 13769 34330 13887 34368
rect 13769 34296 13809 34330
rect 13843 34296 13887 34330
rect 13769 34258 13887 34296
rect 13769 34224 13809 34258
rect 13843 34224 13887 34258
rect 13769 34186 13887 34224
rect 13769 34152 13809 34186
rect 13843 34152 13887 34186
rect 13769 34114 13887 34152
rect 13769 34080 13809 34114
rect 13843 34080 13887 34114
rect 13769 34042 13887 34080
rect 13769 34008 13809 34042
rect 13843 34008 13887 34042
rect 13769 33970 13887 34008
rect 13769 33936 13809 33970
rect 13843 33936 13887 33970
rect 13769 33898 13887 33936
rect 13769 33864 13809 33898
rect 13843 33864 13887 33898
rect 13769 33826 13887 33864
rect 13769 33792 13809 33826
rect 13843 33792 13887 33826
rect 13769 33754 13887 33792
rect 13769 33720 13809 33754
rect 13843 33720 13887 33754
rect 13769 33682 13887 33720
rect 13769 33648 13809 33682
rect 13843 33648 13887 33682
rect 13769 33610 13887 33648
rect 13769 33576 13809 33610
rect 13843 33576 13887 33610
rect 13769 33538 13887 33576
rect 13769 33504 13809 33538
rect 13843 33504 13887 33538
rect 13769 33466 13887 33504
rect 13769 33432 13809 33466
rect 13843 33432 13887 33466
rect 13769 33394 13887 33432
rect 13769 33360 13809 33394
rect 13843 33360 13887 33394
rect 13769 33322 13887 33360
rect 13769 33288 13809 33322
rect 13843 33288 13887 33322
rect 13769 33250 13887 33288
rect 13769 33216 13809 33250
rect 13843 33216 13887 33250
rect 13769 33178 13887 33216
rect 13769 33144 13809 33178
rect 13843 33144 13887 33178
rect 13769 33106 13887 33144
rect 13769 33072 13809 33106
rect 13843 33072 13887 33106
rect 13769 33034 13887 33072
rect 13769 33000 13809 33034
rect 13843 33000 13887 33034
rect 13769 32962 13887 33000
rect 13769 32928 13809 32962
rect 13843 32928 13887 32962
rect 13769 32890 13887 32928
rect 13769 32856 13809 32890
rect 13843 32856 13887 32890
rect 13769 32818 13887 32856
rect 13769 32784 13809 32818
rect 13843 32784 13887 32818
rect 13769 32746 13887 32784
rect 13769 32712 13809 32746
rect 13843 32712 13887 32746
rect 13769 32674 13887 32712
rect 13769 32640 13809 32674
rect 13843 32640 13887 32674
rect 13769 32602 13887 32640
rect 13769 32568 13809 32602
rect 13843 32568 13887 32602
rect 13769 32530 13887 32568
rect 13769 32496 13809 32530
rect 13843 32496 13887 32530
rect 13769 32458 13887 32496
rect 13769 32424 13809 32458
rect 13843 32424 13887 32458
rect 13769 32386 13887 32424
rect 13769 32352 13809 32386
rect 13843 32352 13887 32386
rect 13769 32314 13887 32352
rect 13769 32280 13809 32314
rect 13843 32280 13887 32314
rect 13769 32242 13887 32280
rect 13769 32208 13809 32242
rect 13843 32208 13887 32242
rect 13769 32170 13887 32208
rect 13769 32136 13809 32170
rect 13843 32136 13887 32170
rect 13769 32098 13887 32136
rect 13769 32064 13809 32098
rect 13843 32064 13887 32098
rect 13769 32026 13887 32064
rect 13769 31992 13809 32026
rect 13843 31992 13887 32026
rect 13769 31954 13887 31992
rect 13769 31920 13809 31954
rect 13843 31920 13887 31954
rect 13769 31882 13887 31920
rect 13769 31848 13809 31882
rect 13843 31848 13887 31882
rect 13769 31810 13887 31848
rect 13769 31776 13809 31810
rect 13843 31776 13887 31810
rect 13769 31738 13887 31776
rect 13769 31704 13809 31738
rect 13843 31704 13887 31738
rect 13769 31666 13887 31704
rect 13769 31632 13809 31666
rect 13843 31632 13887 31666
rect 13769 31594 13887 31632
rect 13769 31560 13809 31594
rect 13843 31560 13887 31594
rect 13769 31522 13887 31560
rect 13769 31488 13809 31522
rect 13843 31488 13887 31522
rect 13769 31450 13887 31488
rect 13769 31416 13809 31450
rect 13843 31416 13887 31450
rect 13769 31378 13887 31416
rect 13769 31344 13809 31378
rect 13843 31344 13887 31378
rect 13769 31306 13887 31344
rect 13769 31272 13809 31306
rect 13843 31272 13887 31306
rect 13769 31234 13887 31272
rect 13769 31200 13809 31234
rect 13843 31200 13887 31234
rect 13769 31162 13887 31200
rect 13769 31128 13809 31162
rect 13843 31128 13887 31162
rect 13769 31090 13887 31128
rect 13769 31056 13809 31090
rect 13843 31056 13887 31090
rect 13769 31018 13887 31056
rect 13769 30984 13809 31018
rect 13843 30984 13887 31018
rect 13769 30946 13887 30984
rect 13769 30912 13809 30946
rect 13843 30912 13887 30946
rect 13769 30874 13887 30912
rect 13769 30840 13809 30874
rect 13843 30840 13887 30874
rect 13769 30802 13887 30840
rect 13769 30768 13809 30802
rect 13843 30768 13887 30802
rect 13769 30730 13887 30768
rect 13769 30696 13809 30730
rect 13843 30696 13887 30730
rect 13769 30658 13887 30696
rect 13769 30624 13809 30658
rect 13843 30624 13887 30658
rect 13769 30586 13887 30624
rect 13769 30552 13809 30586
rect 13843 30552 13887 30586
rect 13769 30514 13887 30552
rect 13769 30480 13809 30514
rect 13843 30480 13887 30514
rect 13769 30442 13887 30480
rect 13769 30408 13809 30442
rect 13843 30408 13887 30442
rect 13769 30370 13887 30408
rect 13769 30336 13809 30370
rect 13843 30336 13887 30370
rect 13769 30298 13887 30336
rect 1195 30272 10091 30281
rect 1119 30264 10091 30272
tri 10091 30264 10108 30281 sw
rect 13769 30264 13809 30298
rect 13843 30264 13887 30298
rect 1119 30243 10108 30264
tri 10108 30243 10129 30264 sw
rect 1119 30234 10129 30243
rect 1119 30200 1161 30234
rect 1195 30230 10129 30234
tri 10129 30230 10142 30243 sw
rect 1195 30227 10142 30230
rect 1195 30200 4944 30227
rect 1119 30162 4944 30200
rect 1119 30128 1161 30162
rect 1195 30128 4944 30162
rect 1119 30090 4944 30128
rect 1119 30056 1161 30090
rect 1195 30056 4944 30090
rect 1119 30018 4944 30056
rect 1119 29984 1161 30018
rect 1195 29984 4944 30018
rect 1119 29946 4944 29984
rect 1119 29912 1161 29946
rect 1195 29912 4944 29946
rect 1119 29874 4944 29912
rect 1119 29840 1161 29874
rect 1195 29840 4944 29874
rect 1119 29802 4944 29840
rect 1119 29768 1161 29802
rect 1195 29768 4944 29802
rect 1119 29730 4944 29768
rect 1119 29696 1161 29730
rect 1195 29696 4944 29730
rect 1119 29658 4944 29696
rect 1119 29624 1161 29658
rect 1195 29624 4944 29658
rect 1119 29586 4944 29624
rect 1119 29552 1161 29586
rect 1195 29552 4944 29586
rect 1119 29514 4944 29552
rect 1119 29480 1161 29514
rect 1195 29480 4944 29514
rect 1119 29442 4944 29480
rect 1119 29408 1161 29442
rect 1195 29408 4944 29442
rect 1119 29407 4944 29408
rect 7236 29407 7745 30227
rect 10037 30226 10142 30227
tri 10142 30226 10146 30230 sw
rect 13769 30226 13887 30264
rect 10037 30192 10146 30226
tri 10146 30192 10180 30226 sw
rect 13769 30192 13809 30226
rect 13843 30192 13887 30226
rect 10037 30171 10180 30192
tri 10180 30171 10201 30192 sw
rect 10037 30158 10201 30171
tri 10201 30158 10214 30171 sw
rect 10037 30154 10214 30158
tri 10214 30154 10218 30158 sw
rect 13769 30154 13887 30192
rect 10037 30120 10218 30154
tri 10218 30120 10252 30154 sw
rect 13769 30120 13809 30154
rect 13843 30120 13887 30154
rect 10037 30099 10252 30120
tri 10252 30099 10273 30120 sw
rect 10037 30086 10273 30099
tri 10273 30086 10286 30099 sw
rect 10037 30082 10286 30086
tri 10286 30082 10290 30086 sw
rect 13769 30082 13887 30120
rect 10037 30081 10290 30082
tri 10290 30081 10291 30082 sw
rect 10037 29553 10291 30081
rect 10037 29544 10282 29553
tri 10282 29544 10291 29553 nw
rect 13769 30048 13809 30082
rect 13843 30048 13887 30082
rect 13769 30010 13887 30048
rect 13769 29976 13809 30010
rect 13843 29976 13887 30010
rect 13769 29938 13887 29976
rect 13769 29904 13809 29938
rect 13843 29904 13887 29938
rect 13769 29866 13887 29904
rect 13769 29832 13809 29866
rect 13843 29832 13887 29866
rect 13769 29794 13887 29832
rect 13769 29760 13809 29794
rect 13843 29760 13887 29794
rect 13769 29722 13887 29760
rect 13769 29688 13809 29722
rect 13843 29688 13887 29722
rect 13769 29650 13887 29688
rect 13769 29616 13809 29650
rect 13843 29616 13887 29650
rect 13769 29578 13887 29616
rect 13769 29544 13809 29578
rect 13843 29544 13887 29578
rect 10037 29523 10261 29544
tri 10261 29523 10282 29544 nw
rect 10037 29510 10248 29523
tri 10248 29510 10261 29523 nw
rect 10037 29506 10244 29510
tri 10244 29506 10248 29510 nw
rect 13769 29506 13887 29544
rect 10037 29472 10210 29506
tri 10210 29472 10244 29506 nw
rect 13769 29472 13809 29506
rect 13843 29472 13887 29506
rect 10037 29451 10189 29472
tri 10189 29451 10210 29472 nw
rect 10037 29438 10176 29451
tri 10176 29438 10189 29451 nw
rect 10037 29434 10172 29438
tri 10172 29434 10176 29438 nw
rect 13769 29434 13887 29472
rect 10037 29407 10138 29434
rect 1119 29400 10138 29407
tri 10138 29400 10172 29434 nw
rect 13769 29400 13809 29434
rect 13843 29400 13887 29434
rect 1119 29379 10117 29400
tri 10117 29379 10138 29400 nw
rect 1119 29370 10104 29379
rect 1119 29336 1161 29370
rect 1195 29366 10104 29370
tri 10104 29366 10117 29379 nw
rect 1195 29362 10100 29366
tri 10100 29362 10104 29366 nw
rect 13769 29362 13887 29400
rect 1195 29353 10091 29362
tri 10091 29353 10100 29362 nw
rect 1195 29336 1442 29353
rect 1119 29298 1442 29336
rect 1119 29264 1161 29298
rect 1195 29264 1442 29298
rect 1119 29226 1442 29264
rect 1119 29192 1161 29226
rect 1195 29192 1442 29226
rect 1119 29154 1442 29192
rect 1119 29120 1161 29154
rect 1195 29120 1442 29154
rect 1119 29082 1442 29120
rect 1119 29048 1161 29082
rect 1195 29048 1442 29082
rect 1119 29010 1442 29048
rect 1119 28976 1161 29010
rect 1195 28976 1442 29010
rect 1119 28938 1442 28976
rect 1119 28904 1161 28938
rect 1195 28904 1442 28938
rect 13769 29328 13809 29362
rect 13843 29328 13887 29362
rect 13769 29290 13887 29328
rect 13769 29256 13809 29290
rect 13843 29256 13887 29290
rect 13769 29218 13887 29256
rect 13769 29184 13809 29218
rect 13843 29184 13887 29218
rect 13769 29146 13887 29184
rect 13769 29112 13809 29146
rect 13843 29112 13887 29146
rect 13769 29074 13887 29112
rect 13769 29040 13809 29074
rect 13843 29040 13887 29074
rect 13769 29002 13887 29040
rect 13769 28968 13809 29002
rect 13843 28968 13887 29002
rect 13769 28930 13887 28968
rect 1119 28866 1442 28904
tri 1846 28896 1859 28909 se
rect 1859 28896 13157 28909
tri 13157 28896 13170 28909 sw
rect 13769 28896 13809 28930
rect 13843 28896 13887 28930
tri 1831 28881 1846 28896 se
rect 1846 28881 13170 28896
tri 1825 28875 1831 28881 se
rect 1831 28875 13170 28881
tri 13170 28875 13191 28896 sw
rect 1119 28832 1161 28866
rect 1195 28832 1442 28866
rect 1119 28794 1442 28832
rect 1119 28760 1161 28794
rect 1195 28760 1442 28794
rect 1119 28722 1442 28760
rect 1119 28688 1161 28722
rect 1195 28688 1442 28722
rect 1119 28650 1442 28688
rect 1119 28616 1161 28650
rect 1195 28616 1442 28650
rect 1119 28578 1442 28616
rect 1119 28544 1161 28578
rect 1195 28544 1442 28578
rect 1119 28506 1442 28544
rect 1119 28472 1161 28506
rect 1195 28472 1442 28506
rect 1119 28434 1442 28472
rect 1119 28400 1161 28434
rect 1195 28400 1442 28434
rect 1119 28362 1442 28400
rect 1119 28328 1161 28362
rect 1195 28328 1442 28362
rect 1119 28290 1442 28328
rect 1119 28256 1161 28290
rect 1195 28256 1442 28290
rect 1119 28218 1442 28256
rect 1119 28184 1161 28218
rect 1195 28184 1442 28218
rect 1119 28146 1442 28184
rect 1119 28112 1161 28146
rect 1195 28112 1442 28146
rect 1119 28074 1442 28112
rect 1119 28040 1161 28074
rect 1195 28040 1442 28074
rect 1119 28002 1442 28040
rect 1119 27968 1161 28002
rect 1195 27968 1442 28002
rect 1119 27930 1442 27968
rect 1119 27896 1161 27930
rect 1195 27896 1442 27930
rect 1119 27858 1442 27896
rect 1119 27824 1161 27858
rect 1195 27824 1442 27858
rect 1119 27786 1442 27824
rect 1119 27752 1161 27786
rect 1195 27752 1442 27786
rect 1119 27714 1442 27752
rect 1119 27680 1161 27714
rect 1195 27680 1442 27714
rect 1119 27642 1442 27680
rect 1119 27608 1161 27642
rect 1195 27608 1442 27642
rect 1119 27570 1442 27608
rect 1119 27536 1161 27570
rect 1195 27536 1442 27570
rect 1119 27498 1442 27536
rect 1119 27464 1161 27498
rect 1195 27464 1442 27498
rect 1119 27426 1442 27464
rect 1119 27392 1161 27426
rect 1195 27392 1442 27426
rect 1119 27354 1442 27392
rect 1119 27320 1161 27354
rect 1195 27320 1442 27354
rect 1119 27282 1442 27320
rect 1119 27248 1161 27282
rect 1195 27248 1442 27282
rect 1119 27210 1442 27248
rect 1119 27176 1161 27210
rect 1195 27176 1442 27210
rect 1119 27138 1442 27176
rect 1119 27104 1161 27138
rect 1195 27104 1442 27138
rect 1119 27066 1442 27104
tri 1659 28709 1825 28875 se
rect 1825 28709 1982 28875
rect 1659 28553 1982 28709
rect 13032 28862 13191 28875
tri 13191 28862 13204 28875 sw
rect 13032 28858 13204 28862
tri 13204 28858 13208 28862 sw
rect 13769 28858 13887 28896
rect 13032 28824 13208 28858
tri 13208 28824 13242 28858 sw
rect 13769 28824 13809 28858
rect 13843 28824 13887 28858
rect 13032 28803 13242 28824
tri 13242 28803 13263 28824 sw
rect 13032 28790 13263 28803
tri 13263 28790 13276 28803 sw
rect 13032 28786 13276 28790
tri 13276 28786 13280 28790 sw
rect 13769 28786 13887 28824
rect 13032 28752 13280 28786
tri 13280 28752 13314 28786 sw
rect 13769 28752 13809 28786
rect 13843 28752 13887 28786
rect 13032 28744 13314 28752
tri 13314 28744 13322 28752 sw
rect 13032 28731 13322 28744
tri 13322 28731 13335 28744 sw
rect 13032 28718 13335 28731
tri 13335 28718 13348 28731 sw
rect 13769 28727 13887 28752
rect 14099 34707 14122 34741
rect 14156 34707 14219 34741
rect 14099 34669 14219 34707
rect 14099 34635 14122 34669
rect 14156 34635 14219 34669
rect 14099 34597 14219 34635
rect 14099 34563 14122 34597
rect 14156 34563 14219 34597
rect 14099 34525 14219 34563
rect 14099 34491 14122 34525
rect 14156 34491 14219 34525
rect 14099 34453 14219 34491
rect 14099 34419 14122 34453
rect 14156 34419 14219 34453
rect 14099 34381 14219 34419
rect 14099 34347 14122 34381
rect 14156 34347 14219 34381
rect 14099 34309 14219 34347
rect 14099 34275 14122 34309
rect 14156 34275 14219 34309
rect 14099 34237 14219 34275
rect 14099 34203 14122 34237
rect 14156 34203 14219 34237
rect 14099 34165 14219 34203
rect 14099 34131 14122 34165
rect 14156 34131 14219 34165
rect 14099 34093 14219 34131
rect 14099 34059 14122 34093
rect 14156 34059 14219 34093
rect 14099 34021 14219 34059
rect 14099 33987 14122 34021
rect 14156 33987 14219 34021
rect 14099 33949 14219 33987
rect 14099 33915 14122 33949
rect 14156 33915 14219 33949
rect 14099 33877 14219 33915
rect 14099 33843 14122 33877
rect 14156 33843 14219 33877
rect 14099 33805 14219 33843
rect 14099 33771 14122 33805
rect 14156 33771 14219 33805
rect 14099 33733 14219 33771
rect 14099 33699 14122 33733
rect 14156 33699 14219 33733
rect 14099 33661 14219 33699
rect 14099 33627 14122 33661
rect 14156 33627 14219 33661
rect 14099 33589 14219 33627
rect 14099 33555 14122 33589
rect 14156 33555 14219 33589
rect 14099 33517 14219 33555
rect 14099 33483 14122 33517
rect 14156 33483 14219 33517
rect 14099 33445 14219 33483
rect 14099 33411 14122 33445
rect 14156 33411 14219 33445
rect 14099 33373 14219 33411
rect 14099 33339 14122 33373
rect 14156 33339 14219 33373
rect 14099 33301 14219 33339
rect 14099 33267 14122 33301
rect 14156 33267 14219 33301
rect 14099 33229 14219 33267
rect 14099 33195 14122 33229
rect 14156 33195 14219 33229
rect 14099 33157 14219 33195
rect 14099 33123 14122 33157
rect 14156 33123 14219 33157
rect 14099 33085 14219 33123
rect 14099 33051 14122 33085
rect 14156 33051 14219 33085
rect 14099 33013 14219 33051
rect 14099 32979 14122 33013
rect 14156 32979 14219 33013
rect 14099 32941 14219 32979
rect 14099 32907 14122 32941
rect 14156 32907 14219 32941
rect 14099 32869 14219 32907
rect 14099 32835 14122 32869
rect 14156 32835 14219 32869
rect 14099 32797 14219 32835
rect 14099 32763 14122 32797
rect 14156 32763 14219 32797
rect 14099 32725 14219 32763
rect 14099 32691 14122 32725
rect 14156 32691 14219 32725
rect 14099 32653 14219 32691
rect 14099 32619 14122 32653
rect 14156 32619 14219 32653
rect 14099 32581 14219 32619
rect 14099 32547 14122 32581
rect 14156 32547 14219 32581
rect 14099 32509 14219 32547
rect 14099 32475 14122 32509
rect 14156 32475 14219 32509
rect 14099 32437 14219 32475
rect 14099 32403 14122 32437
rect 14156 32403 14219 32437
rect 14099 32365 14219 32403
rect 14099 32331 14122 32365
rect 14156 32331 14219 32365
rect 14099 32293 14219 32331
rect 14099 32259 14122 32293
rect 14156 32259 14219 32293
rect 14099 32221 14219 32259
rect 14099 32187 14122 32221
rect 14156 32187 14219 32221
rect 14099 32149 14219 32187
rect 14099 32115 14122 32149
rect 14156 32115 14219 32149
rect 14099 32077 14219 32115
rect 14099 32043 14122 32077
rect 14156 32043 14219 32077
rect 14099 32005 14219 32043
rect 14099 31971 14122 32005
rect 14156 31971 14219 32005
rect 14099 31933 14219 31971
rect 14099 31899 14122 31933
rect 14156 31899 14219 31933
rect 14099 31861 14219 31899
rect 14099 31827 14122 31861
rect 14156 31827 14219 31861
rect 14099 31789 14219 31827
rect 14099 31755 14122 31789
rect 14156 31755 14219 31789
rect 14099 31717 14219 31755
rect 14099 31683 14122 31717
rect 14156 31683 14219 31717
rect 14099 31645 14219 31683
rect 14099 31611 14122 31645
rect 14156 31611 14219 31645
rect 14099 31573 14219 31611
rect 14099 31539 14122 31573
rect 14156 31539 14219 31573
rect 14099 31501 14219 31539
rect 14099 31467 14122 31501
rect 14156 31467 14219 31501
rect 14099 31429 14219 31467
rect 14099 31395 14122 31429
rect 14156 31395 14219 31429
rect 14099 31357 14219 31395
rect 14099 31323 14122 31357
rect 14156 31323 14219 31357
rect 14099 31285 14219 31323
rect 14099 31251 14122 31285
rect 14156 31251 14219 31285
rect 14099 31213 14219 31251
rect 14099 31179 14122 31213
rect 14156 31179 14219 31213
rect 14099 31141 14219 31179
rect 14099 31107 14122 31141
rect 14156 31107 14219 31141
rect 14099 31069 14219 31107
rect 14099 31035 14122 31069
rect 14156 31035 14219 31069
rect 14099 30997 14219 31035
rect 14099 30963 14122 30997
rect 14156 30963 14219 30997
rect 14099 30925 14219 30963
rect 14099 30891 14122 30925
rect 14156 30891 14219 30925
rect 14099 30853 14219 30891
rect 14099 30819 14122 30853
rect 14156 30819 14219 30853
rect 14099 30781 14219 30819
rect 14099 30747 14122 30781
rect 14156 30747 14219 30781
rect 14099 30709 14219 30747
rect 14099 30675 14122 30709
rect 14156 30675 14219 30709
rect 14099 30637 14219 30675
rect 14099 30603 14122 30637
rect 14156 30603 14219 30637
rect 14099 30565 14219 30603
rect 14099 30531 14122 30565
rect 14156 30531 14219 30565
rect 14099 30493 14219 30531
rect 14099 30459 14122 30493
rect 14156 30459 14219 30493
rect 14099 30421 14219 30459
rect 14099 30387 14122 30421
rect 14156 30387 14219 30421
rect 14099 30349 14219 30387
rect 14099 30315 14122 30349
rect 14156 30315 14219 30349
rect 14099 30277 14219 30315
rect 14099 30243 14122 30277
rect 14156 30243 14219 30277
rect 14099 30205 14219 30243
rect 14099 30171 14122 30205
rect 14156 30171 14219 30205
rect 14099 30133 14219 30171
rect 14099 30099 14122 30133
rect 14156 30099 14219 30133
rect 14099 30061 14219 30099
rect 14099 30027 14122 30061
rect 14156 30027 14219 30061
rect 14099 29989 14219 30027
rect 14099 29955 14122 29989
rect 14156 29955 14219 29989
rect 14099 29917 14219 29955
rect 14099 29883 14122 29917
rect 14156 29883 14219 29917
rect 14099 29845 14219 29883
rect 14099 29811 14122 29845
rect 14156 29811 14219 29845
rect 14099 29773 14219 29811
rect 14099 29739 14122 29773
rect 14156 29739 14219 29773
rect 14099 29701 14219 29739
rect 14099 29667 14122 29701
rect 14156 29667 14219 29701
rect 14099 29629 14219 29667
rect 14099 29595 14122 29629
rect 14156 29595 14219 29629
rect 14099 29557 14219 29595
rect 14099 29523 14122 29557
rect 14156 29523 14219 29557
rect 14099 29485 14219 29523
rect 14099 29451 14122 29485
rect 14156 29451 14219 29485
rect 14099 29413 14219 29451
rect 14099 29379 14122 29413
rect 14156 29379 14219 29413
rect 14099 29341 14219 29379
rect 14099 29307 14122 29341
rect 14156 29307 14219 29341
rect 14099 29269 14219 29307
rect 14099 29235 14122 29269
rect 14156 29235 14219 29269
rect 14099 29197 14219 29235
rect 14099 29163 14122 29197
rect 14156 29163 14219 29197
rect 14099 29125 14219 29163
rect 14099 29091 14122 29125
rect 14156 29091 14219 29125
rect 14099 29053 14219 29091
rect 14099 29019 14122 29053
rect 14156 29019 14219 29053
rect 14099 28981 14219 29019
rect 14099 28947 14122 28981
rect 14156 28947 14219 28981
rect 14099 28909 14219 28947
rect 14099 28875 14122 28909
rect 14156 28875 14219 28909
rect 14099 28837 14219 28875
rect 14099 28803 14122 28837
rect 14156 28803 14219 28837
rect 14099 28765 14219 28803
rect 14099 28731 14122 28765
rect 14156 28731 14219 28765
rect 13032 28693 13348 28718
tri 13348 28693 13373 28718 sw
rect 14099 28693 14219 28731
rect 13032 28659 13373 28693
tri 13373 28659 13407 28693 sw
rect 14099 28659 14122 28693
rect 14156 28659 14219 28693
rect 13032 28646 13407 28659
tri 13407 28646 13420 28659 sw
rect 13032 28621 13420 28646
tri 13420 28621 13445 28646 sw
rect 14099 28621 14219 28659
rect 13032 28590 13445 28621
tri 13445 28590 13476 28621 sw
rect 13032 28587 13476 28590
tri 13476 28587 13479 28590 sw
rect 14099 28587 14122 28621
rect 14156 28587 14219 28621
rect 13032 28574 13479 28587
tri 13479 28574 13492 28587 sw
rect 13032 28553 13492 28574
rect 1659 28549 13492 28553
tri 13492 28549 13517 28574 sw
rect 14099 28549 14219 28587
rect 1659 28515 13517 28549
tri 13517 28515 13551 28549 sw
rect 14099 28515 14122 28549
rect 14156 28515 14219 28549
rect 1659 28502 2120 28515
tri 2120 28502 2133 28515 nw
tri 12883 28502 12896 28515 ne
rect 12896 28502 13551 28515
tri 13551 28502 13564 28515 sw
rect 1659 28489 2103 28502
rect 1659 27447 1726 28489
rect 1976 28485 2103 28489
tri 2103 28485 2120 28502 nw
tri 12896 28485 12913 28502 ne
rect 12913 28485 13564 28502
rect 1976 28482 2100 28485
tri 2100 28482 2103 28485 nw
tri 12913 28482 12916 28485 ne
rect 12916 28482 13564 28485
rect 1976 27447 2093 28482
tri 2093 28475 2100 28482 nw
tri 12916 28475 12923 28482 ne
tri 2319 28276 2411 28368 se
rect 2411 28335 12604 28368
rect 2411 28276 4939 28335
rect 2319 28219 4939 28276
rect 7231 28219 7750 28335
rect 10042 28276 12604 28335
tri 12604 28276 12696 28368 sw
rect 10042 28219 12696 28276
rect 2319 28168 12696 28219
rect 2509 28022 4482 28048
rect 4481 27906 4482 28022
rect 2509 27880 4482 27906
rect 10500 28022 12473 28048
rect 12472 27906 12473 28022
rect 10500 27880 12473 27906
rect 2320 27719 12696 27764
rect 2320 27652 4939 27719
tri 2320 27552 2420 27652 ne
rect 2420 27603 4939 27652
rect 7231 27603 7750 27719
rect 10042 27652 12696 27719
rect 10042 27603 12596 27652
rect 2420 27552 12596 27603
tri 12596 27552 12696 27652 nw
rect 1659 27440 2093 27447
tri 2093 27440 2104 27451 sw
tri 12912 27440 12923 27451 se
rect 12923 27440 13031 28482
rect 13281 28477 13564 28482
tri 13564 28477 13589 28502 sw
rect 14099 28477 14219 28515
rect 13281 28443 13589 28477
tri 13589 28443 13623 28477 sw
rect 14099 28443 14122 28477
rect 14156 28443 14219 28477
rect 13281 28430 13623 28443
tri 13623 28430 13636 28443 sw
rect 13281 28405 13636 28430
tri 13636 28405 13661 28430 sw
rect 14099 28405 14219 28443
rect 13281 28371 13661 28405
tri 13661 28371 13695 28405 sw
rect 14099 28371 14122 28405
rect 14156 28371 14219 28405
rect 13281 28358 13695 28371
tri 13695 28358 13708 28371 sw
rect 13281 28333 13708 28358
tri 13708 28333 13733 28358 sw
rect 14099 28333 14219 28371
rect 13281 28299 13733 28333
tri 13733 28299 13767 28333 sw
rect 14099 28299 14122 28333
rect 14156 28299 14219 28333
rect 13281 28286 13767 28299
tri 13767 28286 13780 28299 sw
rect 13281 28283 13780 28286
tri 13780 28283 13783 28286 sw
rect 13281 27440 13783 28283
rect 1659 27437 2104 27440
tri 2104 27437 2107 27440 sw
tri 12909 27437 12912 27440 se
rect 12912 27437 13783 27440
rect 1659 27435 2107 27437
tri 2107 27435 2109 27437 sw
tri 12907 27435 12909 27437 se
rect 12909 27435 13783 27437
rect 1659 27422 2109 27435
tri 2109 27422 2122 27435 sw
tri 12894 27422 12907 27435 se
rect 12907 27422 13783 27435
rect 1659 27411 2122 27422
tri 2122 27411 2133 27422 sw
tri 12883 27411 12894 27422 se
rect 12894 27411 13783 27422
rect 1659 27334 13783 27411
rect 1659 27217 1985 27334
tri 1659 27084 1792 27217 ne
rect 1792 27084 1985 27217
rect 13035 27217 13783 27334
rect 13035 27206 13346 27217
tri 13346 27206 13357 27217 nw
rect 13035 27181 13321 27206
tri 13321 27181 13346 27206 nw
rect 13035 27147 13287 27181
tri 13287 27147 13321 27181 nw
rect 13035 27134 13274 27147
tri 13274 27134 13287 27147 nw
rect 13035 27109 13249 27134
tri 13249 27109 13274 27134 nw
rect 13035 27084 13215 27109
tri 1792 27075 1801 27084 ne
rect 1801 27075 13215 27084
tri 13215 27075 13249 27109 nw
rect 1119 27032 1161 27066
rect 1195 27032 1442 27066
tri 1801 27062 1814 27075 ne
rect 1814 27062 13202 27075
tri 13202 27062 13215 27075 nw
tri 1814 27053 1823 27062 ne
rect 1823 27053 13177 27062
tri 1823 27037 1839 27053 ne
rect 1839 27037 13177 27053
tri 13177 27037 13202 27062 nw
rect 1119 26994 1442 27032
tri 1839 27017 1859 27037 ne
rect 1859 27017 13157 27037
tri 13157 27017 13177 27037 nw
rect 1119 26960 1161 26994
rect 1195 26960 1442 26994
rect 1119 26922 1442 26960
rect 1119 26888 1161 26922
rect 1195 26888 1442 26922
rect 1119 26850 1442 26888
rect 1119 26816 1161 26850
rect 1195 26816 1442 26850
rect 1119 26778 1442 26816
rect 1119 26744 1161 26778
rect 1195 26744 1442 26778
rect 1119 26706 1442 26744
rect 1119 26672 1161 26706
rect 1195 26672 1442 26706
rect 1119 26634 1442 26672
rect 1119 26600 1161 26634
rect 1195 26600 1442 26634
rect 1119 26562 1442 26600
rect 1119 26528 1161 26562
rect 1195 26528 1442 26562
rect 1119 26490 1442 26528
rect 1119 26456 1161 26490
rect 1195 26456 1442 26490
rect 1119 26418 1442 26456
rect 1119 26384 1161 26418
rect 1195 26384 1442 26418
rect 1119 26346 1442 26384
rect 1119 26312 1161 26346
rect 1195 26312 1442 26346
rect 1119 26274 1442 26312
rect 1119 26240 1161 26274
rect 1195 26240 1442 26274
rect 1119 26202 1442 26240
rect 1119 26168 1161 26202
rect 1195 26192 1442 26202
rect 1195 26168 1736 26192
rect 1119 26130 1736 26168
rect 1119 26096 1161 26130
rect 1195 26096 1736 26130
rect 1119 26058 1736 26096
rect 1119 26024 1161 26058
rect 1195 26024 1736 26058
tri 2391 26029 2414 26052 se
rect 2414 26029 12578 26052
tri 12578 26029 12601 26052 sw
rect 1119 25986 1736 26024
tri 2357 25995 2391 26029 se
rect 2391 26025 12601 26029
rect 2391 25995 4933 26025
rect 1119 25952 1161 25986
rect 1195 25952 1736 25986
tri 2344 25982 2357 25995 se
rect 2357 25982 4933 25995
rect 1119 25914 1736 25952
rect 1119 25880 1161 25914
rect 1195 25880 1736 25914
tri 2328 25966 2344 25982 se
rect 2344 25966 4933 25982
rect 2328 25909 4933 25966
rect 7225 25909 7757 26025
rect 10049 25995 12601 26025
tri 12601 25995 12635 26029 sw
rect 10049 25982 12635 25995
tri 12635 25982 12648 25995 sw
rect 10049 25966 12648 25982
tri 12648 25966 12664 25982 sw
rect 10049 25909 12664 25966
rect 2328 25880 12664 25909
rect 1119 25842 1736 25880
rect 1119 25808 1161 25842
rect 1195 25808 1736 25842
rect 1119 25770 1736 25808
rect 1119 25736 1161 25770
rect 1195 25736 1736 25770
rect 1119 25698 1736 25736
rect 1119 25664 1161 25698
rect 1195 25664 1736 25698
rect 1119 25626 1736 25664
rect 1119 25592 1161 25626
rect 1195 25592 1736 25626
rect 2528 25759 4472 25781
rect 2528 25643 2546 25759
rect 4454 25643 4472 25759
rect 2528 25621 4472 25643
rect 10510 25759 12454 25781
rect 10510 25643 10528 25759
rect 12436 25643 12454 25759
rect 10510 25621 12454 25643
rect 1119 25554 1736 25592
rect 1119 25520 1161 25554
rect 1195 25520 1736 25554
rect 1119 25482 1736 25520
rect 1119 25448 1161 25482
rect 1195 25448 1736 25482
rect 1119 25410 1736 25448
rect 2326 25493 12662 25520
rect 2326 25428 4933 25493
tri 2326 25419 2335 25428 ne
rect 2335 25419 4933 25428
rect 1119 25376 1161 25410
rect 1195 25376 1736 25410
tri 2335 25406 2348 25419 ne
rect 2348 25406 4933 25419
tri 2348 25381 2373 25406 ne
rect 2373 25381 4933 25406
rect 1119 25338 1736 25376
tri 2373 25348 2406 25381 ne
rect 2406 25377 4933 25381
rect 7225 25377 7757 25493
rect 10049 25428 12662 25493
rect 10049 25419 12653 25428
tri 12653 25419 12662 25428 nw
rect 10049 25406 12640 25419
tri 12640 25406 12653 25419 nw
rect 10049 25381 12615 25406
tri 12615 25381 12640 25406 nw
rect 10049 25377 12582 25381
rect 2406 25348 12582 25377
tri 12582 25348 12615 25381 nw
rect 1119 25304 1161 25338
rect 1195 25304 1736 25338
rect 1119 25266 1736 25304
rect 1119 25232 1161 25266
rect 1195 25232 1736 25266
rect 1119 25202 1736 25232
rect 1119 25194 1237 25202
rect 1119 25160 1161 25194
rect 1195 25160 1237 25194
rect 1119 25122 1237 25160
rect 1119 25088 1161 25122
rect 1195 25088 1237 25122
rect 1119 25050 1237 25088
rect 1119 25016 1161 25050
rect 1195 25016 1237 25050
rect 1119 24978 1237 25016
rect 1119 24944 1161 24978
rect 1195 24944 1237 24978
rect 1119 24906 1237 24944
rect 1119 24872 1161 24906
rect 1195 24872 1237 24906
rect 1119 24834 1237 24872
rect 1119 24800 1161 24834
rect 1195 24800 1237 24834
rect 1119 24762 1237 24800
rect 1119 24728 1161 24762
rect 1195 24728 1237 24762
rect 1119 24690 1237 24728
rect 1119 24656 1161 24690
rect 1195 24656 1237 24690
rect 1119 24618 1237 24656
rect 1119 24584 1161 24618
rect 1195 24584 1237 24618
rect 1119 24546 1237 24584
rect 1119 24512 1161 24546
rect 1195 24512 1237 24546
rect 13527 24543 13783 27217
tri 4890 24542 4891 24543 se
rect 4891 24542 13783 24543
tri 4865 24517 4890 24542 se
rect 4890 24517 13783 24542
rect 1119 24474 1237 24512
tri 4831 24483 4865 24517 se
rect 4865 24489 13783 24517
rect 4865 24483 4945 24489
rect 1119 24440 1161 24474
rect 1195 24440 1237 24474
tri 4818 24470 4831 24483 se
rect 4831 24470 4945 24483
tri 4793 24445 4818 24470 se
rect 4818 24445 4945 24470
rect 1119 24402 1237 24440
tri 4759 24411 4793 24445 se
rect 4793 24411 4945 24445
rect 1119 24368 1161 24402
rect 1195 24368 1237 24402
tri 4746 24398 4759 24411 se
rect 4759 24398 4945 24411
tri 4721 24373 4746 24398 se
rect 4746 24373 4945 24398
rect 1119 24330 1237 24368
rect 1119 24296 1161 24330
rect 1195 24296 1237 24330
rect 1119 24258 1237 24296
rect 1119 24224 1161 24258
rect 1195 24224 1237 24258
rect 1119 24186 1237 24224
rect 1119 24152 1161 24186
rect 1195 24152 1237 24186
rect 1119 24114 1237 24152
rect 1119 24080 1161 24114
rect 1195 24080 1237 24114
rect 1119 24042 1237 24080
rect 1119 24008 1161 24042
rect 1195 24008 1237 24042
rect 1119 23970 1237 24008
rect 1119 23936 1161 23970
rect 1195 23936 1237 23970
rect 1119 23898 1237 23936
rect 1119 23864 1161 23898
rect 1195 23864 1237 23898
rect 1119 23826 1237 23864
rect 1119 23792 1161 23826
rect 1195 23792 1237 23826
tri 4691 24343 4721 24373 se
rect 4721 24343 4945 24373
rect 4691 23815 4945 24343
tri 4691 23797 4709 23815 ne
rect 4709 23797 4945 23815
rect 1119 23754 1237 23792
tri 4709 23763 4743 23797 ne
rect 4743 23763 4945 23797
rect 1119 23720 1161 23754
rect 1195 23720 1237 23754
tri 4743 23750 4756 23763 ne
rect 4756 23750 4945 23763
tri 4756 23725 4781 23750 ne
rect 4781 23725 4945 23750
rect 1119 23682 1237 23720
tri 4781 23691 4815 23725 ne
rect 4815 23691 4945 23725
rect 1119 23648 1161 23682
rect 1195 23648 1237 23682
tri 4815 23678 4828 23691 ne
rect 4828 23678 4945 23691
tri 4828 23653 4853 23678 ne
rect 4853 23669 4945 23678
rect 7237 23669 7744 24489
rect 10036 24041 13783 24489
rect 10036 24038 13780 24041
tri 13780 24038 13783 24041 nw
rect 14099 28261 14219 28299
rect 14099 28227 14122 28261
rect 14156 28227 14219 28261
rect 14099 28189 14219 28227
rect 14099 28155 14122 28189
rect 14156 28155 14219 28189
rect 14099 28117 14219 28155
rect 14099 28083 14122 28117
rect 14156 28083 14219 28117
rect 14099 28045 14219 28083
rect 14099 28011 14122 28045
rect 14156 28011 14219 28045
rect 14099 27973 14219 28011
rect 14099 27939 14122 27973
rect 14156 27939 14219 27973
rect 14099 27901 14219 27939
rect 14099 27867 14122 27901
rect 14156 27867 14219 27901
rect 14099 27829 14219 27867
rect 14099 27795 14122 27829
rect 14156 27795 14219 27829
rect 14099 27757 14219 27795
rect 14099 27723 14122 27757
rect 14156 27723 14219 27757
rect 14099 27685 14219 27723
rect 14099 27651 14122 27685
rect 14156 27651 14219 27685
rect 14099 27613 14219 27651
rect 14099 27579 14122 27613
rect 14156 27579 14219 27613
rect 14099 27541 14219 27579
rect 14099 27507 14122 27541
rect 14156 27507 14219 27541
rect 14099 27469 14219 27507
rect 14099 27435 14122 27469
rect 14156 27435 14219 27469
rect 14099 27397 14219 27435
rect 14099 27363 14122 27397
rect 14156 27363 14219 27397
rect 14099 27325 14219 27363
rect 14099 27291 14122 27325
rect 14156 27291 14219 27325
rect 14099 27253 14219 27291
rect 14099 27219 14122 27253
rect 14156 27219 14219 27253
rect 14099 27181 14219 27219
rect 14099 27147 14122 27181
rect 14156 27147 14219 27181
rect 14099 27109 14219 27147
rect 14099 27075 14122 27109
rect 14156 27075 14219 27109
rect 14099 27037 14219 27075
rect 14099 27003 14122 27037
rect 14156 27003 14219 27037
rect 14099 26965 14219 27003
rect 14099 26931 14122 26965
rect 14156 26931 14219 26965
rect 14099 26893 14219 26931
rect 14099 26859 14122 26893
rect 14156 26859 14219 26893
rect 14099 26821 14219 26859
rect 14099 26787 14122 26821
rect 14156 26787 14219 26821
rect 14099 26749 14219 26787
rect 14099 26715 14122 26749
rect 14156 26715 14219 26749
rect 14099 26677 14219 26715
rect 14099 26643 14122 26677
rect 14156 26643 14219 26677
rect 14099 26605 14219 26643
rect 14099 26571 14122 26605
rect 14156 26571 14219 26605
rect 14099 26533 14219 26571
rect 14099 26499 14122 26533
rect 14156 26499 14219 26533
rect 14099 26461 14219 26499
rect 14099 26427 14122 26461
rect 14156 26427 14219 26461
rect 14099 26389 14219 26427
rect 14099 26355 14122 26389
rect 14156 26355 14219 26389
rect 14099 26317 14219 26355
rect 14099 26283 14122 26317
rect 14156 26283 14219 26317
rect 14099 26245 14219 26283
rect 14099 26211 14122 26245
rect 14156 26211 14219 26245
rect 14099 26173 14219 26211
rect 14099 26139 14122 26173
rect 14156 26139 14219 26173
rect 14099 26101 14219 26139
rect 14099 26067 14122 26101
rect 14156 26067 14219 26101
rect 14099 26029 14219 26067
rect 14099 25995 14122 26029
rect 14156 25995 14219 26029
rect 14099 25957 14219 25995
rect 14099 25923 14122 25957
rect 14156 25923 14219 25957
rect 14099 25885 14219 25923
rect 14099 25851 14122 25885
rect 14156 25851 14219 25885
rect 14099 25813 14219 25851
rect 14099 25779 14122 25813
rect 14156 25779 14219 25813
rect 14099 25741 14219 25779
rect 14099 25707 14122 25741
rect 14156 25707 14219 25741
rect 14099 25669 14219 25707
rect 14099 25635 14122 25669
rect 14156 25635 14219 25669
rect 14099 25597 14219 25635
rect 14099 25563 14122 25597
rect 14156 25563 14219 25597
rect 14099 25525 14219 25563
rect 14099 25491 14122 25525
rect 14156 25491 14219 25525
rect 14099 25453 14219 25491
rect 14099 25419 14122 25453
rect 14156 25419 14219 25453
rect 14099 25381 14219 25419
rect 14099 25347 14122 25381
rect 14156 25347 14219 25381
rect 14099 25309 14219 25347
rect 14099 25275 14122 25309
rect 14156 25275 14219 25309
rect 14099 25237 14219 25275
rect 14099 25203 14122 25237
rect 14156 25203 14219 25237
rect 14099 25165 14219 25203
rect 14099 25131 14122 25165
rect 14156 25131 14219 25165
rect 14099 25093 14219 25131
rect 14099 25059 14122 25093
rect 14156 25059 14219 25093
rect 14099 25021 14219 25059
rect 14099 24987 14122 25021
rect 14156 24987 14219 25021
rect 14099 24949 14219 24987
rect 14099 24915 14122 24949
rect 14156 24915 14219 24949
rect 14099 24877 14219 24915
rect 14099 24843 14122 24877
rect 14156 24843 14219 24877
rect 14099 24805 14219 24843
rect 14099 24771 14122 24805
rect 14156 24771 14219 24805
rect 14099 24733 14219 24771
rect 14099 24699 14122 24733
rect 14156 24699 14219 24733
rect 14099 24661 14219 24699
rect 14099 24627 14122 24661
rect 14156 24627 14219 24661
rect 14099 24589 14219 24627
rect 14099 24555 14122 24589
rect 14156 24555 14219 24589
rect 14099 24517 14219 24555
rect 14099 24483 14122 24517
rect 14156 24483 14219 24517
rect 14099 24445 14219 24483
rect 14099 24411 14122 24445
rect 14156 24411 14219 24445
rect 14099 24373 14219 24411
rect 14099 24339 14122 24373
rect 14156 24339 14219 24373
rect 14099 24301 14219 24339
rect 14099 24267 14122 24301
rect 14156 24267 14219 24301
rect 14099 24229 14219 24267
rect 14099 24195 14122 24229
rect 14156 24195 14219 24229
rect 14099 24157 14219 24195
rect 14099 24123 14122 24157
rect 14156 24123 14219 24157
rect 14099 24085 14219 24123
rect 14099 24051 14122 24085
rect 14156 24051 14219 24085
rect 10036 24013 13755 24038
tri 13755 24013 13780 24038 nw
rect 14099 24013 14219 24051
rect 10036 23979 13721 24013
tri 13721 23979 13755 24013 nw
rect 14099 23979 14122 24013
rect 14156 23979 14219 24013
rect 10036 23966 13708 23979
tri 13708 23966 13721 23979 nw
rect 10036 23941 13683 23966
tri 13683 23941 13708 23966 nw
rect 14099 23941 14219 23979
rect 10036 23907 13649 23941
tri 13649 23907 13683 23941 nw
rect 14099 23907 14122 23941
rect 14156 23907 14219 23941
rect 10036 23894 13636 23907
tri 13636 23894 13649 23907 nw
rect 10036 23869 13611 23894
tri 13611 23869 13636 23894 nw
rect 14099 23869 14219 23907
rect 10036 23835 13577 23869
tri 13577 23835 13611 23869 nw
rect 14099 23835 14122 23869
rect 14156 23835 14219 23869
rect 10036 23822 13564 23835
tri 13564 23822 13577 23835 nw
rect 10036 23797 13539 23822
tri 13539 23797 13564 23822 nw
rect 14099 23797 14219 23835
rect 10036 23763 13505 23797
tri 13505 23763 13539 23797 nw
rect 14099 23763 14122 23797
rect 14156 23763 14219 23797
rect 10036 23750 13492 23763
tri 13492 23750 13505 23763 nw
rect 10036 23725 13467 23750
tri 13467 23725 13492 23750 nw
rect 14099 23725 14219 23763
rect 10036 23691 13433 23725
tri 13433 23691 13467 23725 nw
rect 14099 23691 14122 23725
rect 14156 23691 14219 23725
rect 10036 23678 13420 23691
tri 13420 23678 13433 23691 nw
rect 10036 23669 13395 23678
rect 4853 23653 13395 23669
tri 13395 23653 13420 23678 nw
rect 14099 23653 14219 23691
rect 1119 23610 1237 23648
tri 4853 23619 4887 23653 ne
rect 4887 23619 13361 23653
tri 13361 23619 13395 23653 nw
rect 14099 23619 14122 23653
rect 14156 23619 14219 23653
tri 4887 23615 4891 23619 ne
rect 4891 23615 13357 23619
tri 13357 23615 13361 23619 nw
rect 1119 23576 1161 23610
rect 1195 23576 1237 23610
rect 1119 23538 1237 23576
rect 1119 23504 1161 23538
rect 1195 23504 1237 23538
rect 1119 23466 1237 23504
rect 1119 23432 1161 23466
rect 1195 23432 1237 23466
rect 1119 23394 1237 23432
rect 14099 23581 14219 23619
rect 14099 23547 14122 23581
rect 14156 23547 14219 23581
rect 14099 23509 14219 23547
rect 14099 23475 14122 23509
rect 14156 23475 14219 23509
rect 14099 23437 14219 23475
rect 1119 23360 1161 23394
rect 1195 23360 1237 23394
rect 1119 23322 1237 23360
rect 1119 23288 1161 23322
rect 1195 23288 1237 23322
rect 1119 23250 1237 23288
rect 1119 23216 1161 23250
rect 1195 23216 1237 23250
rect 1119 23178 1237 23216
rect 1119 23144 1161 23178
rect 1195 23144 1237 23178
rect 1119 23106 1237 23144
rect 1119 23072 1161 23106
rect 1195 23072 1237 23106
rect 1119 23034 1237 23072
rect 1119 23000 1161 23034
rect 1195 23000 1237 23034
rect 1119 22962 1237 23000
rect 1119 22928 1161 22962
rect 1195 22928 1237 22962
rect 1119 22890 1237 22928
rect 1119 22856 1161 22890
rect 1195 22856 1237 22890
rect 1119 22818 1237 22856
rect 1119 22784 1161 22818
rect 1195 22784 1237 22818
rect 1119 22746 1237 22784
rect 1119 22712 1161 22746
rect 1195 22712 1237 22746
rect 1119 22674 1237 22712
rect 1119 22640 1161 22674
rect 1195 22640 1237 22674
rect 1119 22602 1237 22640
rect 1119 22568 1161 22602
rect 1195 22568 1237 22602
rect 1119 22530 1237 22568
rect 1119 22496 1161 22530
rect 1195 22496 1237 22530
rect 1119 22458 1237 22496
rect 1119 22424 1161 22458
rect 1195 22424 1237 22458
rect 1119 22386 1237 22424
rect 1119 22352 1161 22386
rect 1195 22352 1237 22386
rect 1119 22314 1237 22352
rect 1119 22280 1161 22314
rect 1195 22280 1237 22314
rect 1119 22242 1237 22280
rect 1119 22208 1161 22242
rect 1195 22208 1237 22242
rect 1119 22170 1237 22208
rect 1119 22136 1161 22170
rect 1195 22136 1237 22170
rect 1119 22098 1237 22136
rect 1119 22064 1161 22098
rect 1195 22064 1237 22098
rect 1119 22026 1237 22064
rect 1119 21992 1161 22026
rect 1195 21992 1237 22026
rect 1119 21954 1237 21992
rect 1119 21920 1161 21954
rect 1195 21920 1237 21954
rect 1119 21882 1237 21920
rect 1119 21848 1161 21882
rect 1195 21848 1237 21882
rect 1119 21810 1237 21848
rect 1119 21776 1161 21810
rect 1195 21776 1237 21810
rect 1119 21738 1237 21776
rect 1119 21704 1161 21738
rect 1195 21704 1237 21738
rect 1119 21666 1237 21704
rect 1119 21632 1161 21666
rect 1195 21632 1237 21666
rect 1119 21594 1237 21632
rect 1119 21560 1161 21594
rect 1195 21560 1237 21594
rect 1119 21522 1237 21560
rect 1119 21488 1161 21522
rect 1195 21488 1237 21522
rect 1119 21450 1237 21488
rect 1119 21416 1161 21450
rect 1195 21416 1237 21450
rect 1119 21378 1237 21416
rect 1119 21344 1161 21378
rect 1195 21344 1237 21378
rect 1119 21306 1237 21344
rect 1119 21272 1161 21306
rect 1195 21272 1237 21306
rect 1119 21234 1237 21272
rect 1119 21200 1161 21234
rect 1195 21200 1237 21234
rect 1119 21162 1237 21200
rect 1119 21128 1161 21162
rect 1195 21128 1237 21162
rect 1119 21090 1237 21128
rect 1119 21056 1161 21090
rect 1195 21056 1237 21090
rect 1119 21018 1237 21056
rect 1119 20984 1161 21018
rect 1195 20984 1237 21018
rect 1119 20946 1237 20984
rect 1119 20912 1161 20946
rect 1195 20912 1237 20946
rect 1119 20874 1237 20912
rect 1119 20840 1161 20874
rect 1195 20840 1237 20874
rect 1119 20802 1237 20840
rect 1119 20768 1161 20802
rect 1195 20768 1237 20802
rect 1119 20730 1237 20768
rect 1119 20696 1161 20730
rect 1195 20696 1237 20730
rect 1119 20658 1237 20696
rect 1119 20624 1161 20658
rect 1195 20624 1237 20658
rect 1119 20586 1237 20624
rect 1119 20552 1161 20586
rect 1195 20552 1237 20586
rect 1119 20514 1237 20552
rect 1119 20480 1161 20514
rect 1195 20480 1237 20514
rect 1119 20442 1237 20480
rect 1119 20408 1161 20442
rect 1195 20408 1237 20442
rect 1119 20370 1237 20408
rect 1119 20336 1161 20370
rect 1195 20336 1237 20370
rect 1119 20298 1237 20336
rect 1119 20264 1161 20298
rect 1195 20264 1237 20298
rect 1119 20226 1237 20264
rect 1119 20192 1161 20226
rect 1195 20192 1237 20226
rect 1119 20154 1237 20192
rect 1119 20120 1161 20154
rect 1195 20120 1237 20154
rect 1119 20082 1237 20120
rect 1119 20048 1161 20082
rect 1195 20048 1237 20082
rect 1119 20010 1237 20048
rect 1119 19976 1161 20010
rect 1195 19976 1237 20010
rect 1119 19938 1237 19976
rect 1119 19904 1161 19938
rect 1195 19904 1237 19938
rect 1119 19866 1237 19904
rect 1119 19832 1161 19866
rect 1195 19832 1237 19866
rect 1119 19794 1237 19832
rect 1119 19760 1161 19794
rect 1195 19760 1237 19794
rect 1119 19722 1237 19760
rect 1119 19688 1161 19722
rect 1195 19688 1237 19722
rect 1119 19650 1237 19688
rect 1119 19616 1161 19650
rect 1195 19616 1237 19650
rect 1119 19578 1237 19616
rect 1119 19544 1161 19578
rect 1195 19544 1237 19578
rect 1119 19506 1237 19544
rect 1119 19472 1161 19506
rect 1195 19472 1237 19506
rect 1119 19434 1237 19472
rect 1119 19400 1161 19434
rect 1195 19400 1237 19434
rect 1119 19362 1237 19400
rect 1119 19328 1161 19362
rect 1195 19328 1237 19362
rect 1119 19290 1237 19328
rect 1119 19256 1161 19290
rect 1195 19256 1237 19290
rect 1119 19218 1237 19256
rect 1119 19184 1161 19218
rect 1195 19184 1237 19218
rect 1119 19146 1237 19184
rect 1119 19112 1161 19146
rect 1195 19112 1237 19146
rect 1119 19074 1237 19112
rect 1119 19040 1161 19074
rect 1195 19040 1237 19074
rect 1119 19002 1237 19040
rect 1119 18968 1161 19002
rect 1195 18968 1237 19002
rect 1119 18930 1237 18968
rect 1119 18896 1161 18930
rect 1195 18896 1237 18930
rect 1119 18858 1237 18896
rect 1119 18824 1161 18858
rect 1195 18824 1237 18858
rect 1119 18786 1237 18824
rect 1119 18752 1161 18786
rect 1195 18752 1237 18786
rect 1119 18714 1237 18752
rect 1119 18680 1161 18714
rect 1195 18680 1237 18714
rect 1119 18642 1237 18680
rect 1119 18608 1161 18642
rect 1195 18608 1237 18642
rect 1119 18570 1237 18608
rect 1119 18536 1161 18570
rect 1195 18536 1237 18570
rect 1119 18498 1237 18536
rect 1119 18464 1161 18498
rect 1195 18464 1237 18498
rect 1119 18426 1237 18464
rect 1119 18392 1161 18426
rect 1195 18392 1237 18426
rect 1119 18354 1237 18392
rect 1119 18320 1161 18354
rect 1195 18320 1237 18354
rect 1119 18282 1237 18320
rect 1119 18248 1161 18282
rect 1195 18248 1237 18282
rect 1119 18210 1237 18248
rect 1119 18176 1161 18210
rect 1195 18176 1237 18210
rect 1119 18138 1237 18176
rect 1119 18104 1161 18138
rect 1195 18104 1237 18138
rect 1119 18066 1237 18104
rect 1119 18032 1161 18066
rect 1195 18032 1237 18066
rect 1119 17994 1237 18032
rect 1119 17960 1161 17994
rect 1195 17960 1237 17994
rect 1119 17922 1237 17960
rect 1119 17888 1161 17922
rect 1195 17888 1237 17922
rect 1119 17850 1237 17888
rect 1119 17816 1161 17850
rect 1195 17816 1237 17850
rect 1119 17778 1237 17816
rect 1119 17744 1161 17778
rect 1195 17744 1237 17778
rect 1119 17706 1237 17744
rect 1119 17672 1161 17706
rect 1195 17672 1237 17706
rect 1119 17634 1237 17672
rect 1119 17600 1161 17634
rect 1195 17600 1237 17634
rect 1119 17562 1237 17600
rect 1119 17528 1161 17562
rect 1195 17528 1237 17562
rect 1119 17490 1237 17528
rect 1119 17456 1161 17490
rect 1195 17456 1237 17490
rect 1119 17418 1237 17456
rect 1119 17384 1161 17418
rect 1195 17384 1237 17418
rect 1119 17346 1237 17384
rect 1119 17312 1161 17346
rect 1195 17312 1237 17346
rect 1119 17274 1237 17312
rect 1119 17240 1161 17274
rect 1195 17240 1237 17274
rect 1119 17202 1237 17240
rect 1119 17168 1161 17202
rect 1195 17168 1237 17202
rect 1119 17130 1237 17168
rect 1119 17096 1161 17130
rect 1195 17096 1237 17130
rect 1119 17058 1237 17096
rect 1119 17024 1161 17058
rect 1195 17024 1237 17058
rect 1119 16986 1237 17024
rect 1119 16952 1161 16986
rect 1195 16952 1237 16986
rect 1119 16914 1237 16952
rect 1119 16880 1161 16914
rect 1195 16880 1237 16914
rect 1119 16842 1237 16880
rect 1119 16808 1161 16842
rect 1195 16808 1237 16842
rect 1119 16770 1237 16808
rect 1119 16736 1161 16770
rect 1195 16736 1237 16770
rect 1119 16698 1237 16736
rect 1119 16664 1161 16698
rect 1195 16664 1237 16698
rect 1119 16626 1237 16664
rect 1119 16592 1161 16626
rect 1195 16592 1237 16626
rect 1119 16554 1237 16592
rect 1119 16520 1161 16554
rect 1195 16520 1237 16554
rect 1119 16482 1237 16520
rect 1119 16448 1161 16482
rect 1195 16448 1237 16482
rect 1119 16410 1237 16448
rect 1119 16376 1161 16410
rect 1195 16376 1237 16410
rect 1119 16338 1237 16376
rect 1119 16304 1161 16338
rect 1195 16304 1237 16338
rect 1119 16266 1237 16304
rect 1119 16232 1161 16266
rect 1195 16232 1237 16266
rect 1119 16194 1237 16232
rect 1119 16160 1161 16194
rect 1195 16160 1237 16194
rect 1119 16122 1237 16160
rect 1119 16088 1161 16122
rect 1195 16088 1237 16122
rect 1119 16050 1237 16088
rect 1119 16016 1161 16050
rect 1195 16016 1237 16050
rect 1119 15978 1237 16016
rect 1119 15944 1161 15978
rect 1195 15944 1237 15978
rect 1119 15906 1237 15944
rect 1119 15872 1161 15906
rect 1195 15872 1237 15906
rect 1119 15834 1237 15872
rect 1119 15800 1161 15834
rect 1195 15800 1237 15834
rect 1119 15762 1237 15800
rect 1119 15728 1161 15762
rect 1195 15728 1237 15762
rect 1119 15690 1237 15728
rect 1119 15656 1161 15690
rect 1195 15656 1237 15690
rect 1119 15618 1237 15656
rect 1119 15584 1161 15618
rect 1195 15584 1237 15618
rect 1119 15546 1237 15584
rect 1119 15512 1161 15546
rect 1195 15512 1237 15546
rect 1119 15474 1237 15512
rect 1119 15440 1161 15474
rect 1195 15440 1237 15474
rect 1119 15402 1237 15440
rect 1119 15368 1161 15402
rect 1195 15368 1237 15402
rect 1119 15319 1237 15368
rect 13769 23397 13888 23428
rect 13769 23363 13809 23397
rect 13843 23363 13888 23397
rect 13769 23325 13888 23363
rect 13769 23291 13809 23325
rect 13843 23291 13888 23325
rect 13769 23253 13888 23291
rect 13769 23219 13809 23253
rect 13843 23219 13888 23253
rect 13769 23181 13888 23219
rect 13769 23147 13809 23181
rect 13843 23147 13888 23181
rect 13769 23109 13888 23147
rect 13769 23075 13809 23109
rect 13843 23075 13888 23109
rect 13769 23037 13888 23075
rect 13769 23003 13809 23037
rect 13843 23003 13888 23037
rect 13769 22965 13888 23003
rect 13769 22931 13809 22965
rect 13843 22931 13888 22965
rect 13769 22893 13888 22931
rect 13769 22859 13809 22893
rect 13843 22859 13888 22893
rect 13769 22821 13888 22859
rect 13769 22787 13809 22821
rect 13843 22787 13888 22821
rect 13769 22749 13888 22787
rect 13769 22715 13809 22749
rect 13843 22715 13888 22749
rect 13769 22677 13888 22715
rect 13769 22643 13809 22677
rect 13843 22643 13888 22677
rect 13769 22605 13888 22643
rect 13769 22571 13809 22605
rect 13843 22571 13888 22605
rect 13769 22533 13888 22571
rect 13769 22499 13809 22533
rect 13843 22499 13888 22533
rect 13769 22461 13888 22499
rect 13769 22427 13809 22461
rect 13843 22427 13888 22461
rect 13769 22389 13888 22427
rect 13769 22355 13809 22389
rect 13843 22355 13888 22389
rect 13769 22317 13888 22355
rect 13769 22283 13809 22317
rect 13843 22283 13888 22317
rect 13769 22245 13888 22283
rect 13769 22211 13809 22245
rect 13843 22211 13888 22245
rect 13769 22173 13888 22211
rect 13769 22139 13809 22173
rect 13843 22139 13888 22173
rect 13769 22101 13888 22139
rect 13769 22067 13809 22101
rect 13843 22067 13888 22101
rect 13769 22029 13888 22067
rect 13769 21995 13809 22029
rect 13843 21995 13888 22029
rect 13769 21957 13888 21995
rect 13769 21923 13809 21957
rect 13843 21923 13888 21957
rect 13769 21885 13888 21923
rect 13769 21851 13809 21885
rect 13843 21851 13888 21885
rect 13769 21813 13888 21851
rect 13769 21779 13809 21813
rect 13843 21779 13888 21813
rect 13769 21741 13888 21779
rect 13769 21707 13809 21741
rect 13843 21707 13888 21741
rect 13769 21669 13888 21707
rect 13769 21635 13809 21669
rect 13843 21635 13888 21669
rect 13769 21597 13888 21635
rect 13769 21563 13809 21597
rect 13843 21563 13888 21597
rect 13769 21525 13888 21563
rect 13769 21491 13809 21525
rect 13843 21491 13888 21525
rect 13769 21453 13888 21491
rect 13769 21419 13809 21453
rect 13843 21419 13888 21453
rect 13769 21381 13888 21419
rect 13769 21347 13809 21381
rect 13843 21347 13888 21381
rect 13769 21309 13888 21347
rect 13769 21275 13809 21309
rect 13843 21275 13888 21309
rect 13769 21237 13888 21275
rect 13769 21203 13809 21237
rect 13843 21203 13888 21237
rect 13769 21165 13888 21203
rect 13769 21131 13809 21165
rect 13843 21131 13888 21165
rect 13769 21093 13888 21131
rect 13769 21059 13809 21093
rect 13843 21059 13888 21093
rect 13769 21021 13888 21059
rect 13769 20987 13809 21021
rect 13843 20987 13888 21021
rect 13769 20949 13888 20987
rect 13769 20915 13809 20949
rect 13843 20915 13888 20949
rect 13769 20877 13888 20915
rect 13769 20843 13809 20877
rect 13843 20843 13888 20877
rect 13769 20805 13888 20843
rect 13769 20771 13809 20805
rect 13843 20771 13888 20805
rect 13769 20733 13888 20771
rect 13769 20699 13809 20733
rect 13843 20699 13888 20733
rect 13769 20661 13888 20699
rect 13769 20627 13809 20661
rect 13843 20627 13888 20661
rect 13769 20589 13888 20627
rect 13769 20555 13809 20589
rect 13843 20555 13888 20589
rect 13769 20517 13888 20555
rect 13769 20483 13809 20517
rect 13843 20483 13888 20517
rect 13769 20445 13888 20483
rect 13769 20411 13809 20445
rect 13843 20411 13888 20445
rect 13769 20373 13888 20411
rect 13769 20339 13809 20373
rect 13843 20339 13888 20373
rect 13769 20301 13888 20339
rect 13769 20267 13809 20301
rect 13843 20267 13888 20301
rect 13769 20229 13888 20267
rect 13769 20195 13809 20229
rect 13843 20195 13888 20229
rect 13769 20157 13888 20195
rect 13769 20123 13809 20157
rect 13843 20123 13888 20157
rect 13769 20085 13888 20123
rect 13769 20051 13809 20085
rect 13843 20051 13888 20085
rect 13769 20013 13888 20051
rect 13769 19979 13809 20013
rect 13843 19979 13888 20013
rect 13769 19941 13888 19979
rect 13769 19907 13809 19941
rect 13843 19907 13888 19941
rect 13769 19869 13888 19907
rect 13769 19835 13809 19869
rect 13843 19835 13888 19869
rect 13769 19797 13888 19835
rect 13769 19763 13809 19797
rect 13843 19763 13888 19797
rect 13769 19725 13888 19763
rect 13769 19691 13809 19725
rect 13843 19691 13888 19725
rect 13769 19653 13888 19691
rect 13769 19619 13809 19653
rect 13843 19619 13888 19653
rect 13769 19581 13888 19619
rect 13769 19547 13809 19581
rect 13843 19547 13888 19581
rect 13769 19509 13888 19547
rect 13769 19475 13809 19509
rect 13843 19475 13888 19509
rect 13769 19437 13888 19475
rect 13769 19403 13809 19437
rect 13843 19403 13888 19437
rect 13769 19365 13888 19403
rect 13769 19331 13809 19365
rect 13843 19331 13888 19365
rect 13769 19293 13888 19331
rect 13769 19259 13809 19293
rect 13843 19259 13888 19293
rect 13769 19221 13888 19259
rect 13769 19187 13809 19221
rect 13843 19187 13888 19221
rect 13769 19149 13888 19187
rect 13769 19115 13809 19149
rect 13843 19115 13888 19149
rect 13769 19077 13888 19115
rect 13769 19043 13809 19077
rect 13843 19043 13888 19077
rect 13769 19005 13888 19043
rect 13769 18971 13809 19005
rect 13843 18971 13888 19005
rect 13769 18933 13888 18971
rect 13769 18899 13809 18933
rect 13843 18899 13888 18933
rect 13769 18861 13888 18899
rect 13769 18827 13809 18861
rect 13843 18827 13888 18861
rect 13769 18789 13888 18827
rect 13769 18755 13809 18789
rect 13843 18755 13888 18789
rect 13769 18717 13888 18755
rect 13769 18683 13809 18717
rect 13843 18683 13888 18717
rect 13769 18645 13888 18683
rect 13769 18611 13809 18645
rect 13843 18611 13888 18645
rect 13769 18573 13888 18611
rect 13769 18539 13809 18573
rect 13843 18539 13888 18573
rect 13769 18501 13888 18539
rect 13769 18467 13809 18501
rect 13843 18467 13888 18501
rect 13769 18429 13888 18467
rect 13769 18395 13809 18429
rect 13843 18395 13888 18429
rect 13769 18357 13888 18395
rect 13769 18323 13809 18357
rect 13843 18323 13888 18357
rect 13769 18285 13888 18323
rect 13769 18251 13809 18285
rect 13843 18251 13888 18285
rect 13769 18213 13888 18251
rect 13769 18179 13809 18213
rect 13843 18179 13888 18213
rect 13769 18141 13888 18179
rect 13769 18107 13809 18141
rect 13843 18107 13888 18141
rect 13769 18069 13888 18107
rect 13769 18035 13809 18069
rect 13843 18035 13888 18069
rect 13769 17997 13888 18035
rect 13769 17963 13809 17997
rect 13843 17963 13888 17997
rect 13769 17925 13888 17963
rect 13769 17891 13809 17925
rect 13843 17891 13888 17925
rect 13769 17853 13888 17891
rect 13769 17819 13809 17853
rect 13843 17819 13888 17853
rect 13769 17781 13888 17819
rect 13769 17747 13809 17781
rect 13843 17747 13888 17781
rect 13769 17709 13888 17747
rect 13769 17675 13809 17709
rect 13843 17675 13888 17709
rect 13769 17637 13888 17675
rect 13769 17603 13809 17637
rect 13843 17603 13888 17637
rect 13769 17565 13888 17603
rect 13769 17531 13809 17565
rect 13843 17531 13888 17565
rect 13769 17493 13888 17531
rect 13769 17459 13809 17493
rect 13843 17459 13888 17493
rect 13769 17421 13888 17459
rect 13769 17387 13809 17421
rect 13843 17387 13888 17421
rect 13769 17349 13888 17387
rect 13769 17315 13809 17349
rect 13843 17315 13888 17349
rect 13769 17277 13888 17315
rect 13769 17243 13809 17277
rect 13843 17243 13888 17277
rect 13769 17205 13888 17243
rect 13769 17171 13809 17205
rect 13843 17171 13888 17205
rect 13769 17133 13888 17171
rect 13769 17099 13809 17133
rect 13843 17099 13888 17133
rect 13769 17061 13888 17099
rect 13769 17027 13809 17061
rect 13843 17027 13888 17061
rect 13769 16989 13888 17027
rect 13769 16955 13809 16989
rect 13843 16955 13888 16989
rect 13769 16917 13888 16955
rect 13769 16883 13809 16917
rect 13843 16883 13888 16917
rect 13769 16845 13888 16883
rect 13769 16811 13809 16845
rect 13843 16811 13888 16845
rect 13769 16773 13888 16811
rect 13769 16739 13809 16773
rect 13843 16739 13888 16773
rect 13769 16701 13888 16739
rect 13769 16667 13809 16701
rect 13843 16667 13888 16701
rect 13769 16629 13888 16667
rect 13769 16595 13809 16629
rect 13843 16595 13888 16629
rect 13769 16557 13888 16595
rect 13769 16523 13809 16557
rect 13843 16523 13888 16557
rect 13769 16485 13888 16523
rect 13769 16451 13809 16485
rect 13843 16451 13888 16485
rect 13769 16413 13888 16451
rect 13769 16379 13809 16413
rect 13843 16379 13888 16413
rect 13769 16341 13888 16379
rect 13769 16307 13809 16341
rect 13843 16307 13888 16341
rect 13769 16269 13888 16307
rect 13769 16235 13809 16269
rect 13843 16235 13888 16269
rect 13769 16197 13888 16235
rect 13769 16163 13809 16197
rect 13843 16163 13888 16197
rect 13769 16125 13888 16163
rect 13769 16091 13809 16125
rect 13843 16091 13888 16125
rect 13769 16053 13888 16091
rect 13769 16019 13809 16053
rect 13843 16019 13888 16053
rect 13769 15981 13888 16019
rect 13769 15947 13809 15981
rect 13843 15947 13888 15981
rect 13769 15909 13888 15947
rect 13769 15875 13809 15909
rect 13843 15875 13888 15909
rect 13769 15837 13888 15875
rect 13769 15803 13809 15837
rect 13843 15803 13888 15837
rect 13769 15765 13888 15803
rect 13769 15731 13809 15765
rect 13843 15731 13888 15765
rect 13769 15693 13888 15731
rect 13769 15659 13809 15693
rect 13843 15659 13888 15693
rect 13769 15621 13888 15659
rect 13769 15587 13809 15621
rect 13843 15587 13888 15621
rect 13769 15549 13888 15587
rect 13769 15515 13809 15549
rect 13843 15515 13888 15549
rect 13769 15477 13888 15515
rect 13769 15443 13809 15477
rect 13843 15443 13888 15477
rect 13769 15405 13888 15443
rect 13769 15371 13809 15405
rect 13843 15371 13888 15405
rect 13769 15319 13888 15371
rect 1119 15278 13888 15319
rect 1119 15244 1298 15278
rect 1332 15244 1370 15278
rect 1404 15244 1442 15278
rect 1476 15244 1514 15278
rect 1548 15244 1586 15278
rect 1620 15244 1658 15278
rect 1692 15244 1730 15278
rect 1764 15244 1802 15278
rect 1836 15244 1874 15278
rect 1908 15244 1946 15278
rect 1980 15244 2018 15278
rect 2052 15244 2090 15278
rect 2124 15244 2162 15278
rect 2196 15244 2234 15278
rect 2268 15244 2306 15278
rect 2340 15244 2378 15278
rect 2412 15244 2450 15278
rect 2484 15244 2522 15278
rect 2556 15244 2594 15278
rect 2628 15244 2666 15278
rect 2700 15244 2738 15278
rect 2772 15244 2810 15278
rect 2844 15244 2882 15278
rect 2916 15244 2954 15278
rect 2988 15244 3026 15278
rect 3060 15244 3098 15278
rect 3132 15244 3170 15278
rect 3204 15244 3242 15278
rect 3276 15244 3314 15278
rect 3348 15244 3386 15278
rect 3420 15244 3458 15278
rect 3492 15244 3530 15278
rect 3564 15244 3602 15278
rect 3636 15244 3674 15278
rect 3708 15244 3746 15278
rect 3780 15244 3818 15278
rect 3852 15244 3890 15278
rect 3924 15244 3962 15278
rect 3996 15244 4034 15278
rect 4068 15244 4106 15278
rect 4140 15244 4178 15278
rect 4212 15244 4250 15278
rect 4284 15244 4322 15278
rect 4356 15244 4394 15278
rect 4428 15244 4466 15278
rect 4500 15244 4538 15278
rect 4572 15244 4610 15278
rect 4644 15244 4682 15278
rect 4716 15244 4754 15278
rect 4788 15244 4826 15278
rect 4860 15244 4898 15278
rect 4932 15244 4970 15278
rect 5004 15244 5042 15278
rect 5076 15244 5114 15278
rect 5148 15244 5186 15278
rect 5220 15244 5258 15278
rect 5292 15244 5330 15278
rect 5364 15244 5402 15278
rect 5436 15244 5474 15278
rect 5508 15244 5546 15278
rect 5580 15244 5618 15278
rect 5652 15244 5690 15278
rect 5724 15244 5762 15278
rect 5796 15244 5834 15278
rect 5868 15244 5906 15278
rect 5940 15244 5978 15278
rect 6012 15244 6050 15278
rect 6084 15244 6122 15278
rect 6156 15244 6194 15278
rect 6228 15244 6266 15278
rect 6300 15244 6338 15278
rect 6372 15244 6410 15278
rect 6444 15244 6482 15278
rect 6516 15244 6554 15278
rect 6588 15244 6626 15278
rect 6660 15244 6698 15278
rect 6732 15244 6770 15278
rect 6804 15244 6842 15278
rect 6876 15244 6914 15278
rect 6948 15244 6986 15278
rect 7020 15244 7058 15278
rect 7092 15244 7130 15278
rect 7164 15244 7202 15278
rect 7236 15244 7274 15278
rect 7308 15244 7346 15278
rect 7380 15244 7418 15278
rect 7452 15244 7490 15278
rect 7524 15244 7562 15278
rect 7596 15244 7634 15278
rect 7668 15244 7706 15278
rect 7740 15244 7778 15278
rect 7812 15244 7850 15278
rect 7884 15244 7922 15278
rect 7956 15244 7994 15278
rect 8028 15244 8066 15278
rect 8100 15244 8138 15278
rect 8172 15244 8210 15278
rect 8244 15244 8282 15278
rect 8316 15244 8354 15278
rect 8388 15244 8426 15278
rect 8460 15244 8498 15278
rect 8532 15244 8570 15278
rect 8604 15244 8642 15278
rect 8676 15244 8714 15278
rect 8748 15244 8786 15278
rect 8820 15244 8858 15278
rect 8892 15244 8930 15278
rect 8964 15244 9002 15278
rect 9036 15244 9074 15278
rect 9108 15244 9146 15278
rect 9180 15244 9218 15278
rect 9252 15244 9290 15278
rect 9324 15244 9362 15278
rect 9396 15244 9434 15278
rect 9468 15244 9506 15278
rect 9540 15244 9578 15278
rect 9612 15244 9650 15278
rect 9684 15244 9722 15278
rect 9756 15244 9794 15278
rect 9828 15244 9866 15278
rect 9900 15244 9938 15278
rect 9972 15244 10010 15278
rect 10044 15244 10082 15278
rect 10116 15244 10154 15278
rect 10188 15244 10226 15278
rect 10260 15244 10298 15278
rect 10332 15244 10370 15278
rect 10404 15244 10442 15278
rect 10476 15244 10514 15278
rect 10548 15244 10586 15278
rect 10620 15244 10658 15278
rect 10692 15244 10730 15278
rect 10764 15244 10802 15278
rect 10836 15244 10874 15278
rect 10908 15244 10946 15278
rect 10980 15244 11018 15278
rect 11052 15244 11090 15278
rect 11124 15244 11162 15278
rect 11196 15244 11234 15278
rect 11268 15244 11306 15278
rect 11340 15244 11378 15278
rect 11412 15244 11450 15278
rect 11484 15244 11522 15278
rect 11556 15244 11594 15278
rect 11628 15244 11666 15278
rect 11700 15244 11738 15278
rect 11772 15244 11810 15278
rect 11844 15244 11882 15278
rect 11916 15244 11954 15278
rect 11988 15244 12026 15278
rect 12060 15244 12098 15278
rect 12132 15244 12170 15278
rect 12204 15244 12242 15278
rect 12276 15244 12314 15278
rect 12348 15244 12386 15278
rect 12420 15244 12458 15278
rect 12492 15244 12530 15278
rect 12564 15244 12602 15278
rect 12636 15244 12674 15278
rect 12708 15244 12746 15278
rect 12780 15244 12818 15278
rect 12852 15244 12890 15278
rect 12924 15244 12962 15278
rect 12996 15244 13034 15278
rect 13068 15244 13106 15278
rect 13140 15244 13178 15278
rect 13212 15244 13250 15278
rect 13284 15244 13322 15278
rect 13356 15244 13394 15278
rect 13428 15244 13466 15278
rect 13500 15244 13538 15278
rect 13572 15244 13610 15278
rect 13644 15244 13682 15278
rect 13716 15244 13888 15278
rect 1119 15201 13888 15244
rect 14099 23403 14122 23437
rect 14156 23403 14219 23437
rect 14099 23365 14219 23403
rect 14099 23331 14122 23365
rect 14156 23331 14219 23365
rect 14099 23293 14219 23331
rect 14099 23259 14122 23293
rect 14156 23259 14219 23293
rect 14099 23221 14219 23259
rect 14099 23187 14122 23221
rect 14156 23187 14219 23221
rect 14099 23149 14219 23187
rect 14099 23115 14122 23149
rect 14156 23115 14219 23149
rect 14099 23077 14219 23115
rect 14099 23043 14122 23077
rect 14156 23043 14219 23077
rect 14099 23005 14219 23043
rect 14099 22971 14122 23005
rect 14156 22971 14219 23005
rect 14099 22933 14219 22971
rect 14099 22899 14122 22933
rect 14156 22899 14219 22933
rect 14099 22861 14219 22899
rect 14099 22827 14122 22861
rect 14156 22827 14219 22861
rect 14099 22789 14219 22827
rect 14099 22755 14122 22789
rect 14156 22755 14219 22789
rect 14099 22717 14219 22755
rect 14099 22683 14122 22717
rect 14156 22683 14219 22717
rect 14099 22645 14219 22683
rect 14099 22611 14122 22645
rect 14156 22611 14219 22645
rect 14099 22573 14219 22611
rect 14099 22539 14122 22573
rect 14156 22539 14219 22573
rect 14099 22501 14219 22539
rect 14099 22467 14122 22501
rect 14156 22467 14219 22501
rect 14099 22429 14219 22467
rect 14099 22395 14122 22429
rect 14156 22395 14219 22429
rect 14099 22357 14219 22395
rect 14099 22323 14122 22357
rect 14156 22323 14219 22357
rect 14099 22285 14219 22323
rect 14099 22251 14122 22285
rect 14156 22251 14219 22285
rect 14099 22213 14219 22251
rect 14099 22179 14122 22213
rect 14156 22179 14219 22213
rect 14099 22141 14219 22179
rect 14099 22107 14122 22141
rect 14156 22107 14219 22141
rect 14099 22069 14219 22107
rect 14099 22035 14122 22069
rect 14156 22035 14219 22069
rect 14099 21997 14219 22035
rect 14099 21963 14122 21997
rect 14156 21963 14219 21997
rect 14099 21925 14219 21963
rect 14099 21891 14122 21925
rect 14156 21891 14219 21925
rect 14099 21853 14219 21891
rect 14099 21819 14122 21853
rect 14156 21819 14219 21853
rect 14099 21781 14219 21819
rect 14099 21747 14122 21781
rect 14156 21747 14219 21781
rect 14099 21709 14219 21747
rect 14099 21675 14122 21709
rect 14156 21675 14219 21709
rect 14099 21637 14219 21675
rect 14099 21603 14122 21637
rect 14156 21603 14219 21637
rect 14099 21565 14219 21603
rect 14099 21531 14122 21565
rect 14156 21531 14219 21565
rect 14099 21493 14219 21531
rect 14099 21459 14122 21493
rect 14156 21459 14219 21493
rect 14099 21421 14219 21459
rect 14099 21387 14122 21421
rect 14156 21387 14219 21421
rect 14099 21349 14219 21387
rect 14099 21315 14122 21349
rect 14156 21315 14219 21349
rect 14099 21277 14219 21315
rect 14099 21243 14122 21277
rect 14156 21243 14219 21277
rect 14099 21205 14219 21243
rect 14099 21171 14122 21205
rect 14156 21171 14219 21205
rect 14099 21133 14219 21171
rect 14099 21099 14122 21133
rect 14156 21099 14219 21133
rect 14099 21061 14219 21099
rect 14099 21027 14122 21061
rect 14156 21027 14219 21061
rect 14099 20989 14219 21027
rect 14099 20955 14122 20989
rect 14156 20955 14219 20989
rect 14099 20917 14219 20955
rect 14099 20883 14122 20917
rect 14156 20883 14219 20917
rect 14099 20845 14219 20883
rect 14099 20811 14122 20845
rect 14156 20811 14219 20845
rect 14099 20773 14219 20811
rect 14099 20739 14122 20773
rect 14156 20739 14219 20773
rect 14099 20701 14219 20739
rect 14099 20667 14122 20701
rect 14156 20667 14219 20701
rect 14099 20629 14219 20667
rect 14099 20595 14122 20629
rect 14156 20595 14219 20629
rect 14099 20557 14219 20595
rect 14099 20523 14122 20557
rect 14156 20523 14219 20557
rect 14099 20485 14219 20523
rect 14099 20451 14122 20485
rect 14156 20451 14219 20485
rect 14099 20413 14219 20451
rect 14099 20379 14122 20413
rect 14156 20379 14219 20413
rect 14099 20341 14219 20379
rect 14099 20307 14122 20341
rect 14156 20307 14219 20341
rect 14099 20269 14219 20307
rect 14099 20235 14122 20269
rect 14156 20235 14219 20269
rect 14099 20197 14219 20235
rect 14099 20163 14122 20197
rect 14156 20163 14219 20197
rect 14099 20125 14219 20163
rect 14099 20091 14122 20125
rect 14156 20091 14219 20125
rect 14099 20053 14219 20091
rect 14099 20019 14122 20053
rect 14156 20019 14219 20053
rect 14099 19981 14219 20019
rect 14099 19947 14122 19981
rect 14156 19947 14219 19981
rect 14099 19909 14219 19947
rect 14099 19875 14122 19909
rect 14156 19875 14219 19909
rect 14099 19837 14219 19875
rect 14099 19803 14122 19837
rect 14156 19803 14219 19837
rect 14099 19765 14219 19803
rect 14099 19731 14122 19765
rect 14156 19731 14219 19765
rect 14099 19693 14219 19731
rect 14099 19659 14122 19693
rect 14156 19659 14219 19693
rect 14099 19621 14219 19659
rect 14099 19587 14122 19621
rect 14156 19587 14219 19621
rect 14099 19549 14219 19587
rect 14099 19515 14122 19549
rect 14156 19515 14219 19549
rect 14099 19477 14219 19515
rect 14099 19443 14122 19477
rect 14156 19443 14219 19477
rect 14099 19405 14219 19443
rect 14099 19371 14122 19405
rect 14156 19371 14219 19405
rect 14099 19333 14219 19371
rect 14099 19299 14122 19333
rect 14156 19299 14219 19333
rect 14099 19261 14219 19299
rect 14099 19227 14122 19261
rect 14156 19227 14219 19261
rect 14099 19189 14219 19227
rect 14099 19155 14122 19189
rect 14156 19155 14219 19189
rect 14099 19117 14219 19155
rect 14099 19083 14122 19117
rect 14156 19083 14219 19117
rect 14099 19045 14219 19083
rect 14099 19011 14122 19045
rect 14156 19011 14219 19045
rect 14099 18973 14219 19011
rect 14099 18939 14122 18973
rect 14156 18939 14219 18973
rect 14099 18901 14219 18939
rect 14099 18867 14122 18901
rect 14156 18867 14219 18901
rect 14099 18829 14219 18867
rect 14099 18795 14122 18829
rect 14156 18795 14219 18829
rect 14099 18757 14219 18795
rect 14099 18723 14122 18757
rect 14156 18723 14219 18757
rect 14099 18685 14219 18723
rect 14099 18651 14122 18685
rect 14156 18651 14219 18685
rect 14099 18613 14219 18651
rect 14099 18579 14122 18613
rect 14156 18579 14219 18613
rect 14099 18541 14219 18579
rect 14099 18507 14122 18541
rect 14156 18507 14219 18541
rect 14099 18469 14219 18507
rect 14099 18435 14122 18469
rect 14156 18435 14219 18469
rect 14099 18397 14219 18435
rect 14099 18363 14122 18397
rect 14156 18363 14219 18397
rect 14099 18325 14219 18363
rect 14099 18291 14122 18325
rect 14156 18291 14219 18325
rect 14099 18253 14219 18291
rect 14099 18219 14122 18253
rect 14156 18219 14219 18253
rect 14099 18181 14219 18219
rect 14099 18147 14122 18181
rect 14156 18147 14219 18181
rect 14099 18109 14219 18147
rect 14099 18075 14122 18109
rect 14156 18075 14219 18109
rect 14099 18037 14219 18075
rect 14099 18003 14122 18037
rect 14156 18003 14219 18037
rect 14099 17965 14219 18003
rect 14099 17931 14122 17965
rect 14156 17931 14219 17965
rect 14099 17893 14219 17931
rect 14099 17859 14122 17893
rect 14156 17859 14219 17893
rect 14099 17821 14219 17859
rect 14099 17787 14122 17821
rect 14156 17787 14219 17821
rect 14099 17749 14219 17787
rect 14099 17715 14122 17749
rect 14156 17715 14219 17749
rect 14099 17677 14219 17715
rect 14099 17643 14122 17677
rect 14156 17643 14219 17677
rect 14099 17605 14219 17643
rect 14099 17571 14122 17605
rect 14156 17571 14219 17605
rect 14099 17533 14219 17571
rect 14099 17499 14122 17533
rect 14156 17499 14219 17533
rect 14099 17461 14219 17499
rect 14099 17427 14122 17461
rect 14156 17427 14219 17461
rect 14099 17389 14219 17427
rect 14099 17355 14122 17389
rect 14156 17355 14219 17389
rect 14099 17317 14219 17355
rect 14099 17283 14122 17317
rect 14156 17283 14219 17317
rect 14099 17245 14219 17283
rect 14099 17211 14122 17245
rect 14156 17211 14219 17245
rect 14099 17173 14219 17211
rect 14099 17139 14122 17173
rect 14156 17139 14219 17173
rect 14099 17101 14219 17139
rect 14099 17067 14122 17101
rect 14156 17067 14219 17101
rect 14099 17029 14219 17067
rect 14099 16995 14122 17029
rect 14156 16995 14219 17029
rect 14099 16957 14219 16995
rect 14099 16923 14122 16957
rect 14156 16923 14219 16957
rect 14099 16885 14219 16923
rect 14099 16851 14122 16885
rect 14156 16851 14219 16885
rect 14099 16813 14219 16851
rect 14099 16779 14122 16813
rect 14156 16779 14219 16813
rect 14099 16741 14219 16779
rect 14099 16707 14122 16741
rect 14156 16707 14219 16741
rect 14099 16669 14219 16707
rect 14099 16635 14122 16669
rect 14156 16635 14219 16669
rect 14099 16597 14219 16635
rect 14099 16563 14122 16597
rect 14156 16563 14219 16597
rect 14099 16525 14219 16563
rect 14099 16491 14122 16525
rect 14156 16491 14219 16525
rect 14099 16453 14219 16491
rect 14099 16419 14122 16453
rect 14156 16419 14219 16453
rect 14099 16381 14219 16419
rect 14099 16347 14122 16381
rect 14156 16347 14219 16381
rect 14099 16309 14219 16347
rect 14099 16275 14122 16309
rect 14156 16275 14219 16309
rect 14099 16237 14219 16275
rect 14099 16203 14122 16237
rect 14156 16203 14219 16237
rect 14099 16165 14219 16203
rect 14099 16131 14122 16165
rect 14156 16131 14219 16165
rect 14099 16093 14219 16131
rect 14099 16059 14122 16093
rect 14156 16059 14219 16093
rect 14099 16021 14219 16059
rect 14099 15987 14122 16021
rect 14156 15987 14219 16021
rect 14099 15949 14219 15987
rect 14099 15915 14122 15949
rect 14156 15915 14219 15949
rect 14099 15877 14219 15915
rect 14099 15843 14122 15877
rect 14156 15843 14219 15877
rect 14099 15805 14219 15843
rect 14099 15771 14122 15805
rect 14156 15771 14219 15805
rect 14099 15733 14219 15771
rect 14099 15699 14122 15733
rect 14156 15699 14219 15733
rect 14099 15661 14219 15699
rect 14099 15627 14122 15661
rect 14156 15627 14219 15661
rect 14099 15589 14219 15627
rect 14099 15555 14122 15589
rect 14156 15555 14219 15589
rect 14099 15517 14219 15555
rect 14099 15483 14122 15517
rect 14156 15483 14219 15517
rect 14099 15445 14219 15483
rect 14099 15411 14122 15445
rect 14156 15411 14219 15445
rect 14099 15373 14219 15411
rect 14099 15339 14122 15373
rect 14156 15339 14219 15373
rect 14099 15301 14219 15339
rect 14099 15267 14122 15301
rect 14156 15267 14219 15301
rect 14099 15229 14219 15267
rect 757 15130 807 15164
rect 841 15130 877 15164
rect 757 15092 877 15130
rect 757 15058 807 15092
rect 841 15058 877 15092
rect 757 14966 877 15058
rect 14099 15195 14122 15229
rect 14156 15195 14219 15229
rect 14099 15157 14219 15195
rect 14099 15123 14122 15157
rect 14156 15123 14219 15157
rect 14099 15085 14219 15123
rect 14099 15051 14122 15085
rect 14156 15051 14219 15085
tri 877 14966 914 15003 sw
tri 14062 14966 14099 15003 se
rect 14099 14966 14219 15051
rect 757 14963 914 14966
tri 914 14963 917 14966 sw
tri 14059 14963 14062 14966 se
rect 14062 14963 14219 14966
rect 757 14943 14219 14963
tri 757 14942 758 14943 ne
rect 758 14942 14208 14943
rect 245 14897 430 14935
tri 758 14908 792 14942 ne
rect 792 14908 891 14942
rect 925 14908 963 14942
rect 997 14908 1035 14942
rect 1069 14908 1107 14942
rect 1141 14908 1179 14942
rect 1213 14908 1251 14942
rect 1285 14908 1323 14942
rect 1357 14908 1395 14942
rect 1429 14908 1467 14942
rect 1501 14908 1539 14942
rect 1573 14908 1611 14942
rect 1645 14908 1683 14942
rect 1717 14908 1755 14942
rect 1789 14908 1827 14942
rect 1861 14908 1899 14942
rect 1933 14908 1971 14942
rect 2005 14908 2043 14942
rect 2077 14908 2115 14942
rect 2149 14908 2187 14942
rect 2221 14908 2259 14942
rect 2293 14908 2331 14942
rect 2365 14908 2403 14942
rect 2437 14908 2475 14942
rect 2509 14908 2547 14942
rect 2581 14908 2619 14942
rect 2653 14908 2691 14942
rect 2725 14908 2763 14942
rect 2797 14908 2835 14942
rect 2869 14908 2907 14942
rect 2941 14908 2979 14942
rect 3013 14908 3051 14942
rect 3085 14908 3123 14942
rect 3157 14908 3195 14942
rect 3229 14908 3267 14942
rect 3301 14908 3339 14942
rect 3373 14908 3411 14942
rect 3445 14908 3483 14942
rect 3517 14908 3555 14942
rect 3589 14908 3627 14942
rect 3661 14908 3699 14942
rect 3733 14908 3771 14942
rect 3805 14908 3843 14942
rect 3877 14908 3915 14942
rect 3949 14908 3987 14942
rect 4021 14908 4059 14942
rect 4093 14908 4131 14942
rect 4165 14908 4203 14942
rect 4237 14908 4275 14942
rect 4309 14908 4347 14942
rect 4381 14908 4419 14942
rect 4453 14908 4491 14942
rect 4525 14908 4563 14942
rect 4597 14908 4635 14942
rect 4669 14908 4707 14942
rect 4741 14908 4779 14942
rect 4813 14908 4851 14942
rect 4885 14908 4923 14942
rect 4957 14908 4995 14942
rect 5029 14908 5067 14942
rect 5101 14908 5139 14942
rect 5173 14908 5211 14942
rect 5245 14908 5283 14942
rect 5317 14908 5355 14942
rect 5389 14908 5427 14942
rect 5461 14908 5499 14942
rect 5533 14908 5571 14942
rect 5605 14908 5643 14942
rect 5677 14908 5715 14942
rect 5749 14908 5787 14942
rect 5821 14908 5859 14942
rect 5893 14908 5931 14942
rect 5965 14908 6003 14942
rect 6037 14908 6075 14942
rect 6109 14908 6147 14942
rect 6181 14908 6219 14942
rect 6253 14908 6291 14942
rect 6325 14908 6363 14942
rect 6397 14908 6435 14942
rect 6469 14908 6507 14942
rect 6541 14908 6579 14942
rect 6613 14908 6651 14942
rect 6685 14908 6723 14942
rect 6757 14908 6795 14942
rect 6829 14908 6867 14942
rect 6901 14908 6939 14942
rect 6973 14908 7011 14942
rect 7045 14908 7083 14942
rect 7117 14908 7155 14942
rect 7189 14908 7227 14942
rect 7261 14908 7299 14942
rect 7333 14908 7371 14942
rect 7405 14908 7443 14942
rect 7477 14908 7515 14942
rect 7549 14908 7587 14942
rect 7621 14908 7659 14942
rect 7693 14908 7731 14942
rect 7765 14908 7803 14942
rect 7837 14908 7875 14942
rect 7909 14908 7947 14942
rect 7981 14908 8019 14942
rect 8053 14908 8091 14942
rect 8125 14908 8163 14942
rect 8197 14908 8235 14942
rect 8269 14908 8307 14942
rect 8341 14908 8379 14942
rect 8413 14908 8451 14942
rect 8485 14908 8523 14942
rect 8557 14908 8595 14942
rect 8629 14908 8667 14942
rect 8701 14908 8739 14942
rect 8773 14908 8811 14942
rect 8845 14908 8883 14942
rect 8917 14908 8955 14942
rect 8989 14908 9027 14942
rect 9061 14908 9099 14942
rect 9133 14908 9171 14942
rect 9205 14908 9243 14942
rect 9277 14908 9315 14942
rect 9349 14908 9387 14942
rect 9421 14908 9459 14942
rect 9493 14908 9531 14942
rect 9565 14908 9603 14942
rect 9637 14908 9675 14942
rect 9709 14908 9747 14942
rect 9781 14908 9819 14942
rect 9853 14908 9891 14942
rect 9925 14908 9963 14942
rect 9997 14908 10035 14942
rect 10069 14908 10107 14942
rect 10141 14908 10179 14942
rect 10213 14908 10251 14942
rect 10285 14908 10323 14942
rect 10357 14908 10395 14942
rect 10429 14908 10467 14942
rect 10501 14908 10539 14942
rect 10573 14908 10611 14942
rect 10645 14908 10683 14942
rect 10717 14908 10755 14942
rect 10789 14908 10827 14942
rect 10861 14908 10899 14942
rect 10933 14908 10971 14942
rect 11005 14908 11043 14942
rect 11077 14908 11115 14942
rect 11149 14908 11187 14942
rect 11221 14908 11259 14942
rect 11293 14908 11331 14942
rect 11365 14908 11403 14942
rect 11437 14908 11475 14942
rect 11509 14908 11547 14942
rect 11581 14908 11619 14942
rect 11653 14908 11691 14942
rect 11725 14908 11763 14942
rect 11797 14908 11835 14942
rect 11869 14908 11907 14942
rect 11941 14908 11979 14942
rect 12013 14908 12051 14942
rect 12085 14908 12123 14942
rect 12157 14908 12195 14942
rect 12229 14908 12267 14942
rect 12301 14908 12339 14942
rect 12373 14908 12411 14942
rect 12445 14908 12483 14942
rect 12517 14908 12555 14942
rect 12589 14908 12627 14942
rect 12661 14908 12699 14942
rect 12733 14908 12771 14942
rect 12805 14908 12843 14942
rect 12877 14908 12915 14942
rect 12949 14908 12987 14942
rect 13021 14908 13059 14942
rect 13093 14908 13131 14942
rect 13165 14908 13203 14942
rect 13237 14908 13275 14942
rect 13309 14908 13347 14942
rect 13381 14908 13419 14942
rect 13453 14908 13491 14942
rect 13525 14908 13563 14942
rect 13597 14908 13635 14942
rect 13669 14908 13707 14942
rect 13741 14908 13779 14942
rect 13813 14908 13851 14942
rect 13885 14908 13923 14942
rect 13957 14908 13995 14942
rect 14029 14932 14208 14942
tri 14208 14932 14219 14943 nw
rect 14539 35918 14724 35956
rect 14539 35884 14614 35918
rect 14648 35884 14724 35918
rect 14539 35846 14724 35884
rect 14539 35812 14614 35846
rect 14648 35812 14724 35846
rect 14539 35774 14724 35812
rect 14539 35740 14614 35774
rect 14648 35740 14724 35774
rect 14539 35702 14724 35740
rect 14539 35668 14614 35702
rect 14648 35668 14724 35702
rect 14539 35630 14724 35668
rect 14539 35596 14614 35630
rect 14648 35596 14724 35630
rect 14539 35558 14724 35596
rect 14539 35524 14614 35558
rect 14648 35524 14724 35558
rect 14539 35486 14724 35524
rect 14539 35452 14614 35486
rect 14648 35452 14724 35486
rect 14539 35414 14724 35452
rect 14539 35380 14614 35414
rect 14648 35380 14724 35414
rect 14539 35342 14724 35380
rect 14539 35308 14614 35342
rect 14648 35308 14724 35342
rect 14539 35270 14724 35308
rect 14539 35236 14614 35270
rect 14648 35236 14724 35270
rect 14539 35198 14724 35236
rect 14539 35164 14614 35198
rect 14648 35164 14724 35198
rect 14539 35126 14724 35164
rect 14539 35092 14614 35126
rect 14648 35092 14724 35126
rect 14539 35054 14724 35092
rect 14539 35020 14614 35054
rect 14648 35020 14724 35054
rect 14539 34982 14724 35020
rect 14539 34948 14614 34982
rect 14648 34948 14724 34982
rect 14539 34910 14724 34948
rect 14539 34876 14614 34910
rect 14648 34876 14724 34910
rect 14539 34838 14724 34876
rect 14539 34804 14614 34838
rect 14648 34804 14724 34838
rect 14539 34766 14724 34804
rect 14539 34732 14614 34766
rect 14648 34732 14724 34766
rect 14539 34694 14724 34732
rect 14539 34660 14614 34694
rect 14648 34660 14724 34694
rect 14539 34622 14724 34660
rect 14539 34588 14614 34622
rect 14648 34588 14724 34622
rect 14539 34550 14724 34588
rect 14539 34516 14614 34550
rect 14648 34516 14724 34550
rect 14539 34478 14724 34516
rect 14539 34444 14614 34478
rect 14648 34444 14724 34478
rect 14539 34406 14724 34444
rect 14539 34372 14614 34406
rect 14648 34372 14724 34406
rect 14539 34334 14724 34372
rect 14539 34300 14614 34334
rect 14648 34300 14724 34334
rect 14539 34262 14724 34300
rect 14539 34228 14614 34262
rect 14648 34228 14724 34262
rect 14539 34190 14724 34228
rect 14539 34156 14614 34190
rect 14648 34156 14724 34190
rect 14539 34118 14724 34156
rect 14539 34084 14614 34118
rect 14648 34084 14724 34118
rect 14539 34046 14724 34084
rect 14539 34012 14614 34046
rect 14648 34012 14724 34046
rect 14539 33974 14724 34012
rect 14539 33940 14614 33974
rect 14648 33940 14724 33974
rect 14539 33902 14724 33940
rect 14539 33868 14614 33902
rect 14648 33868 14724 33902
rect 14539 33830 14724 33868
rect 14539 33796 14614 33830
rect 14648 33796 14724 33830
rect 14539 33758 14724 33796
rect 14539 33724 14614 33758
rect 14648 33724 14724 33758
rect 14539 33686 14724 33724
rect 14539 33652 14614 33686
rect 14648 33652 14724 33686
rect 14539 33614 14724 33652
rect 14539 33580 14614 33614
rect 14648 33580 14724 33614
rect 14539 33542 14724 33580
rect 14539 33508 14614 33542
rect 14648 33508 14724 33542
rect 14539 33470 14724 33508
rect 14539 33436 14614 33470
rect 14648 33436 14724 33470
rect 14539 33398 14724 33436
rect 14539 33364 14614 33398
rect 14648 33364 14724 33398
rect 14539 33326 14724 33364
rect 14539 33292 14614 33326
rect 14648 33292 14724 33326
rect 14539 33254 14724 33292
rect 14539 33220 14614 33254
rect 14648 33220 14724 33254
rect 14539 33182 14724 33220
rect 14539 33148 14614 33182
rect 14648 33148 14724 33182
rect 14539 33110 14724 33148
rect 14539 33076 14614 33110
rect 14648 33076 14724 33110
rect 14539 33038 14724 33076
rect 14539 33004 14614 33038
rect 14648 33004 14724 33038
rect 14539 32966 14724 33004
rect 14539 32932 14614 32966
rect 14648 32932 14724 32966
rect 14539 32894 14724 32932
rect 14539 32860 14614 32894
rect 14648 32860 14724 32894
rect 14539 32822 14724 32860
rect 14539 32788 14614 32822
rect 14648 32788 14724 32822
rect 14539 32750 14724 32788
rect 14539 32716 14614 32750
rect 14648 32716 14724 32750
rect 14539 32678 14724 32716
rect 14539 32644 14614 32678
rect 14648 32644 14724 32678
rect 14539 32606 14724 32644
rect 14539 32572 14614 32606
rect 14648 32572 14724 32606
rect 14539 32534 14724 32572
rect 14539 32500 14614 32534
rect 14648 32500 14724 32534
rect 14539 32462 14724 32500
rect 14539 32428 14614 32462
rect 14648 32428 14724 32462
rect 14539 32390 14724 32428
rect 14539 32356 14614 32390
rect 14648 32356 14724 32390
rect 14539 32318 14724 32356
rect 14539 32284 14614 32318
rect 14648 32284 14724 32318
rect 14539 32246 14724 32284
rect 14539 32212 14614 32246
rect 14648 32212 14724 32246
rect 14539 32174 14724 32212
rect 14539 32140 14614 32174
rect 14648 32140 14724 32174
rect 14539 32102 14724 32140
rect 14539 32068 14614 32102
rect 14648 32068 14724 32102
rect 14539 32030 14724 32068
rect 14539 31996 14614 32030
rect 14648 31996 14724 32030
rect 14539 31958 14724 31996
rect 14539 31924 14614 31958
rect 14648 31924 14724 31958
rect 14539 31886 14724 31924
rect 14539 31852 14614 31886
rect 14648 31852 14724 31886
rect 14539 31814 14724 31852
rect 14539 31780 14614 31814
rect 14648 31780 14724 31814
rect 14539 31742 14724 31780
rect 14539 31708 14614 31742
rect 14648 31708 14724 31742
rect 14539 31670 14724 31708
rect 14539 31636 14614 31670
rect 14648 31636 14724 31670
rect 14539 31598 14724 31636
rect 14539 31564 14614 31598
rect 14648 31564 14724 31598
rect 14539 31526 14724 31564
rect 14539 31492 14614 31526
rect 14648 31492 14724 31526
rect 14539 31454 14724 31492
rect 14539 31420 14614 31454
rect 14648 31420 14724 31454
rect 14539 31382 14724 31420
rect 14539 31348 14614 31382
rect 14648 31348 14724 31382
rect 14539 31310 14724 31348
rect 14539 31276 14614 31310
rect 14648 31276 14724 31310
rect 14539 31238 14724 31276
rect 14539 31204 14614 31238
rect 14648 31204 14724 31238
rect 14539 31166 14724 31204
rect 14539 31132 14614 31166
rect 14648 31132 14724 31166
rect 14539 31094 14724 31132
rect 14539 31060 14614 31094
rect 14648 31060 14724 31094
rect 14539 31022 14724 31060
rect 14539 30988 14614 31022
rect 14648 30988 14724 31022
rect 14539 30950 14724 30988
rect 14539 30916 14614 30950
rect 14648 30916 14724 30950
rect 14539 30878 14724 30916
rect 14539 30844 14614 30878
rect 14648 30844 14724 30878
rect 14539 30806 14724 30844
rect 14539 30772 14614 30806
rect 14648 30772 14724 30806
rect 14539 30734 14724 30772
rect 14539 30700 14614 30734
rect 14648 30700 14724 30734
rect 14539 30662 14724 30700
rect 14539 30628 14614 30662
rect 14648 30628 14724 30662
rect 14539 30590 14724 30628
rect 14539 30556 14614 30590
rect 14648 30556 14724 30590
rect 14539 30518 14724 30556
rect 14539 30484 14614 30518
rect 14648 30484 14724 30518
rect 14539 30446 14724 30484
rect 14539 30412 14614 30446
rect 14648 30412 14724 30446
rect 14539 30374 14724 30412
rect 14539 30340 14614 30374
rect 14648 30340 14724 30374
rect 14539 30302 14724 30340
rect 14539 30268 14614 30302
rect 14648 30268 14724 30302
rect 14539 30230 14724 30268
rect 14539 30196 14614 30230
rect 14648 30196 14724 30230
rect 14539 30158 14724 30196
rect 14539 30124 14614 30158
rect 14648 30124 14724 30158
rect 14539 30086 14724 30124
rect 14539 30052 14614 30086
rect 14648 30052 14724 30086
rect 14539 30014 14724 30052
rect 14539 29980 14614 30014
rect 14648 29980 14724 30014
rect 14539 29942 14724 29980
rect 14539 29908 14614 29942
rect 14648 29908 14724 29942
rect 14539 29870 14724 29908
rect 14539 29836 14614 29870
rect 14648 29836 14724 29870
rect 14539 29798 14724 29836
rect 14539 29764 14614 29798
rect 14648 29764 14724 29798
rect 14539 29726 14724 29764
rect 14539 29692 14614 29726
rect 14648 29692 14724 29726
rect 14539 29654 14724 29692
rect 14539 29620 14614 29654
rect 14648 29620 14724 29654
rect 14539 29582 14724 29620
rect 14539 29548 14614 29582
rect 14648 29548 14724 29582
rect 14539 29510 14724 29548
rect 14539 29476 14614 29510
rect 14648 29476 14724 29510
rect 14539 29438 14724 29476
rect 14539 29404 14614 29438
rect 14648 29404 14724 29438
rect 14539 29366 14724 29404
rect 14539 29332 14614 29366
rect 14648 29332 14724 29366
rect 14539 29294 14724 29332
rect 14539 29260 14614 29294
rect 14648 29260 14724 29294
rect 14539 29222 14724 29260
rect 14539 29188 14614 29222
rect 14648 29188 14724 29222
rect 14539 29150 14724 29188
rect 14539 29116 14614 29150
rect 14648 29116 14724 29150
rect 14539 29078 14724 29116
rect 14539 29044 14614 29078
rect 14648 29044 14724 29078
rect 14539 29006 14724 29044
rect 14539 28972 14614 29006
rect 14648 28972 14724 29006
rect 14539 28934 14724 28972
rect 14539 28900 14614 28934
rect 14648 28900 14724 28934
rect 14539 28862 14724 28900
rect 14539 28828 14614 28862
rect 14648 28828 14724 28862
rect 14539 28790 14724 28828
rect 14539 28756 14614 28790
rect 14648 28756 14724 28790
rect 14539 28718 14724 28756
rect 14539 28684 14614 28718
rect 14648 28684 14724 28718
rect 14539 28646 14724 28684
rect 14539 28612 14614 28646
rect 14648 28612 14724 28646
rect 14539 28574 14724 28612
rect 14539 28540 14614 28574
rect 14648 28540 14724 28574
rect 14539 28502 14724 28540
rect 14539 28468 14614 28502
rect 14648 28468 14724 28502
rect 14539 28430 14724 28468
rect 14539 28396 14614 28430
rect 14648 28396 14724 28430
rect 14539 28358 14724 28396
rect 14539 28324 14614 28358
rect 14648 28324 14724 28358
rect 14539 28286 14724 28324
rect 14539 28252 14614 28286
rect 14648 28252 14724 28286
rect 14539 28214 14724 28252
rect 14539 28180 14614 28214
rect 14648 28180 14724 28214
rect 14539 28142 14724 28180
rect 14539 28108 14614 28142
rect 14648 28108 14724 28142
rect 14539 28070 14724 28108
rect 14539 28036 14614 28070
rect 14648 28036 14724 28070
rect 14539 27998 14724 28036
rect 14539 27964 14614 27998
rect 14648 27964 14724 27998
rect 14539 27926 14724 27964
rect 14539 27892 14614 27926
rect 14648 27892 14724 27926
rect 14539 27854 14724 27892
rect 14539 27820 14614 27854
rect 14648 27820 14724 27854
rect 14539 27782 14724 27820
rect 14539 27748 14614 27782
rect 14648 27748 14724 27782
rect 14539 27710 14724 27748
rect 14539 27676 14614 27710
rect 14648 27676 14724 27710
rect 14539 27638 14724 27676
rect 14539 27604 14614 27638
rect 14648 27604 14724 27638
rect 14539 27566 14724 27604
rect 14539 27532 14614 27566
rect 14648 27532 14724 27566
rect 14539 27494 14724 27532
rect 14539 27460 14614 27494
rect 14648 27460 14724 27494
rect 14539 27422 14724 27460
rect 14539 27388 14614 27422
rect 14648 27388 14724 27422
rect 14539 27350 14724 27388
rect 14539 27316 14614 27350
rect 14648 27316 14724 27350
rect 14539 27278 14724 27316
rect 14539 27244 14614 27278
rect 14648 27244 14724 27278
rect 14539 27206 14724 27244
rect 14539 27172 14614 27206
rect 14648 27172 14724 27206
rect 14539 27134 14724 27172
rect 14539 27100 14614 27134
rect 14648 27100 14724 27134
rect 14539 27062 14724 27100
rect 14539 27028 14614 27062
rect 14648 27028 14724 27062
rect 14539 26990 14724 27028
rect 14539 26956 14614 26990
rect 14648 26956 14724 26990
rect 14539 26918 14724 26956
rect 14539 26884 14614 26918
rect 14648 26884 14724 26918
rect 14539 26846 14724 26884
rect 14539 26812 14614 26846
rect 14648 26812 14724 26846
rect 14539 26774 14724 26812
rect 14539 26740 14614 26774
rect 14648 26740 14724 26774
rect 14539 26702 14724 26740
rect 14539 26668 14614 26702
rect 14648 26668 14724 26702
rect 14539 26630 14724 26668
rect 14539 26596 14614 26630
rect 14648 26596 14724 26630
rect 14539 26558 14724 26596
rect 14539 26524 14614 26558
rect 14648 26524 14724 26558
rect 14539 26486 14724 26524
rect 14539 26452 14614 26486
rect 14648 26452 14724 26486
rect 14539 26414 14724 26452
rect 14539 26380 14614 26414
rect 14648 26380 14724 26414
rect 14539 26342 14724 26380
rect 14539 26308 14614 26342
rect 14648 26308 14724 26342
rect 14539 26270 14724 26308
rect 14539 26236 14614 26270
rect 14648 26236 14724 26270
rect 14539 26198 14724 26236
rect 14539 26164 14614 26198
rect 14648 26164 14724 26198
rect 14539 26126 14724 26164
rect 14539 26092 14614 26126
rect 14648 26092 14724 26126
rect 14539 26054 14724 26092
rect 14539 26020 14614 26054
rect 14648 26020 14724 26054
rect 14539 25982 14724 26020
rect 14539 25948 14614 25982
rect 14648 25948 14724 25982
rect 14539 25910 14724 25948
rect 14539 25876 14614 25910
rect 14648 25876 14724 25910
rect 14539 25838 14724 25876
rect 14539 25804 14614 25838
rect 14648 25804 14724 25838
rect 14539 25766 14724 25804
rect 14539 25732 14614 25766
rect 14648 25732 14724 25766
rect 14539 25694 14724 25732
rect 14539 25660 14614 25694
rect 14648 25660 14724 25694
rect 14539 25622 14724 25660
rect 14539 25588 14614 25622
rect 14648 25588 14724 25622
rect 14539 25550 14724 25588
rect 14539 25516 14614 25550
rect 14648 25516 14724 25550
rect 14539 25478 14724 25516
rect 14539 25444 14614 25478
rect 14648 25444 14724 25478
rect 14539 25406 14724 25444
rect 14539 25372 14614 25406
rect 14648 25372 14724 25406
rect 14539 25334 14724 25372
rect 14539 25300 14614 25334
rect 14648 25300 14724 25334
rect 14539 25262 14724 25300
rect 14539 25228 14614 25262
rect 14648 25228 14724 25262
rect 14539 25190 14724 25228
rect 14539 25156 14614 25190
rect 14648 25156 14724 25190
rect 14539 25118 14724 25156
rect 14539 25084 14614 25118
rect 14648 25084 14724 25118
rect 14539 25046 14724 25084
rect 14539 25012 14614 25046
rect 14648 25012 14724 25046
rect 14539 24974 14724 25012
rect 14539 24940 14614 24974
rect 14648 24940 14724 24974
rect 14539 24902 14724 24940
rect 14539 24868 14614 24902
rect 14648 24868 14724 24902
rect 14539 24830 14724 24868
rect 14539 24796 14614 24830
rect 14648 24796 14724 24830
rect 14539 24758 14724 24796
rect 14539 24724 14614 24758
rect 14648 24724 14724 24758
rect 14539 24686 14724 24724
rect 14539 24652 14614 24686
rect 14648 24652 14724 24686
rect 14539 24614 14724 24652
rect 14539 24580 14614 24614
rect 14648 24580 14724 24614
rect 14539 24542 14724 24580
rect 14539 24508 14614 24542
rect 14648 24508 14724 24542
rect 14539 24470 14724 24508
rect 14539 24436 14614 24470
rect 14648 24436 14724 24470
rect 14539 24398 14724 24436
rect 14539 24364 14614 24398
rect 14648 24364 14724 24398
rect 14539 24326 14724 24364
rect 14539 24292 14614 24326
rect 14648 24292 14724 24326
rect 14539 24254 14724 24292
rect 14539 24220 14614 24254
rect 14648 24220 14724 24254
rect 14539 24182 14724 24220
rect 14539 24148 14614 24182
rect 14648 24148 14724 24182
rect 14539 24110 14724 24148
rect 14539 24076 14614 24110
rect 14648 24076 14724 24110
rect 14539 24038 14724 24076
rect 14539 24004 14614 24038
rect 14648 24004 14724 24038
rect 14539 23966 14724 24004
rect 14539 23932 14614 23966
rect 14648 23932 14724 23966
rect 14539 23894 14724 23932
rect 14539 23860 14614 23894
rect 14648 23860 14724 23894
rect 14539 23822 14724 23860
rect 14539 23788 14614 23822
rect 14648 23788 14724 23822
rect 14539 23750 14724 23788
rect 14539 23716 14614 23750
rect 14648 23716 14724 23750
rect 14539 23678 14724 23716
rect 14539 23644 14614 23678
rect 14648 23644 14724 23678
rect 14539 23606 14724 23644
rect 14539 23572 14614 23606
rect 14648 23572 14724 23606
rect 14539 23534 14724 23572
rect 14539 23500 14614 23534
rect 14648 23500 14724 23534
rect 14539 23462 14724 23500
rect 14539 23428 14614 23462
rect 14648 23428 14724 23462
rect 14539 23390 14724 23428
rect 14539 23356 14614 23390
rect 14648 23356 14724 23390
rect 14539 23318 14724 23356
rect 14539 23284 14614 23318
rect 14648 23284 14724 23318
rect 14539 23246 14724 23284
rect 14539 23212 14614 23246
rect 14648 23212 14724 23246
rect 14539 23174 14724 23212
rect 14539 23140 14614 23174
rect 14648 23140 14724 23174
rect 14539 23102 14724 23140
rect 14539 23068 14614 23102
rect 14648 23068 14724 23102
rect 14539 23030 14724 23068
rect 14539 22996 14614 23030
rect 14648 22996 14724 23030
rect 14539 22958 14724 22996
rect 14539 22924 14614 22958
rect 14648 22924 14724 22958
rect 14539 22886 14724 22924
rect 14539 22852 14614 22886
rect 14648 22852 14724 22886
rect 14539 22814 14724 22852
rect 14539 22780 14614 22814
rect 14648 22780 14724 22814
rect 14539 22742 14724 22780
rect 14539 22708 14614 22742
rect 14648 22708 14724 22742
rect 14539 22670 14724 22708
rect 14539 22636 14614 22670
rect 14648 22636 14724 22670
rect 14539 22598 14724 22636
rect 14539 22564 14614 22598
rect 14648 22564 14724 22598
rect 14539 22526 14724 22564
rect 14539 22492 14614 22526
rect 14648 22492 14724 22526
rect 14539 22454 14724 22492
rect 14539 22420 14614 22454
rect 14648 22420 14724 22454
rect 14539 22382 14724 22420
rect 14539 22348 14614 22382
rect 14648 22348 14724 22382
rect 14539 22310 14724 22348
rect 14539 22276 14614 22310
rect 14648 22276 14724 22310
rect 14539 22238 14724 22276
rect 14539 22204 14614 22238
rect 14648 22204 14724 22238
rect 14539 22166 14724 22204
rect 14539 22132 14614 22166
rect 14648 22132 14724 22166
rect 14539 22094 14724 22132
rect 14539 22060 14614 22094
rect 14648 22060 14724 22094
rect 14539 22022 14724 22060
rect 14539 21988 14614 22022
rect 14648 21988 14724 22022
rect 14539 21950 14724 21988
rect 14539 21916 14614 21950
rect 14648 21916 14724 21950
rect 14539 21878 14724 21916
rect 14539 21844 14614 21878
rect 14648 21844 14724 21878
rect 14539 21806 14724 21844
rect 14539 21772 14614 21806
rect 14648 21772 14724 21806
rect 14539 21734 14724 21772
rect 14539 21700 14614 21734
rect 14648 21700 14724 21734
rect 14539 21662 14724 21700
rect 14539 21628 14614 21662
rect 14648 21628 14724 21662
rect 14539 21590 14724 21628
rect 14539 21556 14614 21590
rect 14648 21556 14724 21590
rect 14539 21518 14724 21556
rect 14539 21484 14614 21518
rect 14648 21484 14724 21518
rect 14539 21446 14724 21484
rect 14539 21412 14614 21446
rect 14648 21412 14724 21446
rect 14539 21374 14724 21412
rect 14539 21340 14614 21374
rect 14648 21340 14724 21374
rect 14539 21302 14724 21340
rect 14539 21268 14614 21302
rect 14648 21268 14724 21302
rect 14539 21230 14724 21268
rect 14539 21196 14614 21230
rect 14648 21196 14724 21230
rect 14539 21158 14724 21196
rect 14539 21124 14614 21158
rect 14648 21124 14724 21158
rect 14539 21086 14724 21124
rect 14539 21052 14614 21086
rect 14648 21052 14724 21086
rect 14539 21014 14724 21052
rect 14539 20980 14614 21014
rect 14648 20980 14724 21014
rect 14539 20942 14724 20980
rect 14539 20908 14614 20942
rect 14648 20908 14724 20942
rect 14539 20870 14724 20908
rect 14539 20836 14614 20870
rect 14648 20836 14724 20870
rect 14539 20798 14724 20836
rect 14539 20764 14614 20798
rect 14648 20764 14724 20798
rect 14539 20726 14724 20764
rect 14539 20692 14614 20726
rect 14648 20692 14724 20726
rect 14539 20654 14724 20692
rect 14539 20620 14614 20654
rect 14648 20620 14724 20654
rect 14539 20582 14724 20620
rect 14539 20548 14614 20582
rect 14648 20548 14724 20582
rect 14539 20510 14724 20548
rect 14539 20476 14614 20510
rect 14648 20476 14724 20510
rect 14539 20438 14724 20476
rect 14539 20404 14614 20438
rect 14648 20404 14724 20438
rect 14539 20366 14724 20404
rect 14539 20332 14614 20366
rect 14648 20332 14724 20366
rect 14539 20294 14724 20332
rect 14539 20260 14614 20294
rect 14648 20260 14724 20294
rect 14539 20222 14724 20260
rect 14539 20188 14614 20222
rect 14648 20188 14724 20222
rect 14539 20150 14724 20188
rect 14539 20116 14614 20150
rect 14648 20116 14724 20150
rect 14539 20078 14724 20116
rect 14539 20044 14614 20078
rect 14648 20044 14724 20078
rect 14539 20006 14724 20044
rect 14539 19972 14614 20006
rect 14648 19972 14724 20006
rect 14539 19934 14724 19972
rect 14539 19900 14614 19934
rect 14648 19900 14724 19934
rect 14539 19862 14724 19900
rect 14539 19828 14614 19862
rect 14648 19828 14724 19862
rect 14539 19790 14724 19828
rect 14539 19756 14614 19790
rect 14648 19756 14724 19790
rect 14539 19718 14724 19756
rect 14539 19684 14614 19718
rect 14648 19684 14724 19718
rect 14539 19646 14724 19684
rect 14539 19612 14614 19646
rect 14648 19612 14724 19646
rect 14539 19574 14724 19612
rect 14539 19540 14614 19574
rect 14648 19540 14724 19574
rect 14539 19502 14724 19540
rect 14539 19468 14614 19502
rect 14648 19468 14724 19502
rect 14539 19430 14724 19468
rect 14539 19396 14614 19430
rect 14648 19396 14724 19430
rect 14539 19358 14724 19396
rect 14539 19324 14614 19358
rect 14648 19324 14724 19358
rect 14539 19286 14724 19324
rect 14539 19252 14614 19286
rect 14648 19252 14724 19286
rect 14539 19214 14724 19252
rect 14539 19180 14614 19214
rect 14648 19180 14724 19214
rect 14539 19142 14724 19180
rect 14539 19108 14614 19142
rect 14648 19108 14724 19142
rect 14539 19070 14724 19108
rect 14539 19036 14614 19070
rect 14648 19036 14724 19070
rect 14539 18998 14724 19036
rect 14539 18964 14614 18998
rect 14648 18964 14724 18998
rect 14539 18926 14724 18964
rect 14539 18892 14614 18926
rect 14648 18892 14724 18926
rect 14539 18854 14724 18892
rect 14539 18820 14614 18854
rect 14648 18820 14724 18854
rect 14539 18782 14724 18820
rect 14539 18748 14614 18782
rect 14648 18748 14724 18782
rect 14539 18710 14724 18748
rect 14539 18676 14614 18710
rect 14648 18676 14724 18710
rect 14539 18638 14724 18676
rect 14539 18604 14614 18638
rect 14648 18604 14724 18638
rect 14539 18566 14724 18604
rect 14539 18532 14614 18566
rect 14648 18532 14724 18566
rect 14539 18494 14724 18532
rect 14539 18460 14614 18494
rect 14648 18460 14724 18494
rect 14539 18422 14724 18460
rect 14539 18388 14614 18422
rect 14648 18388 14724 18422
rect 14539 18350 14724 18388
rect 14539 18316 14614 18350
rect 14648 18316 14724 18350
rect 14539 18278 14724 18316
rect 14539 18244 14614 18278
rect 14648 18244 14724 18278
rect 14539 18206 14724 18244
rect 14539 18172 14614 18206
rect 14648 18172 14724 18206
rect 14539 18134 14724 18172
rect 14539 18100 14614 18134
rect 14648 18100 14724 18134
rect 14539 18062 14724 18100
rect 14539 18028 14614 18062
rect 14648 18028 14724 18062
rect 14539 17990 14724 18028
rect 14539 17956 14614 17990
rect 14648 17956 14724 17990
rect 14539 17918 14724 17956
rect 14539 17884 14614 17918
rect 14648 17884 14724 17918
rect 14539 17846 14724 17884
rect 14539 17812 14614 17846
rect 14648 17812 14724 17846
rect 14539 17774 14724 17812
rect 14539 17740 14614 17774
rect 14648 17740 14724 17774
rect 14539 17702 14724 17740
rect 14539 17668 14614 17702
rect 14648 17668 14724 17702
rect 14539 17630 14724 17668
rect 14539 17596 14614 17630
rect 14648 17596 14724 17630
rect 14539 17558 14724 17596
rect 14539 17524 14614 17558
rect 14648 17524 14724 17558
rect 14539 17486 14724 17524
rect 14539 17452 14614 17486
rect 14648 17452 14724 17486
rect 14539 17414 14724 17452
rect 14539 17380 14614 17414
rect 14648 17380 14724 17414
rect 14539 17342 14724 17380
rect 14539 17308 14614 17342
rect 14648 17308 14724 17342
rect 14539 17270 14724 17308
rect 14539 17236 14614 17270
rect 14648 17236 14724 17270
rect 14539 17198 14724 17236
rect 14539 17164 14614 17198
rect 14648 17164 14724 17198
rect 14539 17126 14724 17164
rect 14539 17092 14614 17126
rect 14648 17092 14724 17126
rect 14539 17054 14724 17092
rect 14539 17020 14614 17054
rect 14648 17020 14724 17054
rect 14539 16982 14724 17020
rect 14539 16948 14614 16982
rect 14648 16948 14724 16982
rect 14539 16910 14724 16948
rect 14539 16876 14614 16910
rect 14648 16876 14724 16910
rect 14539 16838 14724 16876
rect 14539 16804 14614 16838
rect 14648 16804 14724 16838
rect 14539 16766 14724 16804
rect 14539 16732 14614 16766
rect 14648 16732 14724 16766
rect 14539 16694 14724 16732
rect 14539 16660 14614 16694
rect 14648 16660 14724 16694
rect 14539 16622 14724 16660
rect 14539 16588 14614 16622
rect 14648 16588 14724 16622
rect 14539 16550 14724 16588
rect 14539 16516 14614 16550
rect 14648 16516 14724 16550
rect 14539 16478 14724 16516
rect 14539 16444 14614 16478
rect 14648 16444 14724 16478
rect 14539 16406 14724 16444
rect 14539 16372 14614 16406
rect 14648 16372 14724 16406
rect 14539 16334 14724 16372
rect 14539 16300 14614 16334
rect 14648 16300 14724 16334
rect 14539 16262 14724 16300
rect 14539 16228 14614 16262
rect 14648 16228 14724 16262
rect 14539 16190 14724 16228
rect 14539 16156 14614 16190
rect 14648 16156 14724 16190
rect 14539 16118 14724 16156
rect 14539 16084 14614 16118
rect 14648 16084 14724 16118
rect 14539 16046 14724 16084
rect 14539 16012 14614 16046
rect 14648 16012 14724 16046
rect 14539 15974 14724 16012
rect 14539 15940 14614 15974
rect 14648 15940 14724 15974
rect 14539 15902 14724 15940
rect 14539 15868 14614 15902
rect 14648 15868 14724 15902
rect 14539 15830 14724 15868
rect 14539 15796 14614 15830
rect 14648 15796 14724 15830
rect 14539 15758 14724 15796
rect 14539 15724 14614 15758
rect 14648 15724 14724 15758
rect 14539 15686 14724 15724
rect 14539 15652 14614 15686
rect 14648 15652 14724 15686
rect 14539 15614 14724 15652
rect 14539 15580 14614 15614
rect 14648 15580 14724 15614
rect 14539 15542 14724 15580
rect 14539 15508 14614 15542
rect 14648 15508 14724 15542
rect 14539 15470 14724 15508
rect 14539 15436 14614 15470
rect 14648 15436 14724 15470
rect 14539 15398 14724 15436
rect 14539 15364 14614 15398
rect 14648 15364 14724 15398
rect 14539 15326 14724 15364
rect 14539 15292 14614 15326
rect 14648 15292 14724 15326
rect 14539 15254 14724 15292
rect 14539 15220 14614 15254
rect 14648 15220 14724 15254
rect 14539 15182 14724 15220
rect 14539 15148 14614 15182
rect 14648 15148 14724 15182
rect 14539 15110 14724 15148
rect 14539 15076 14614 15110
rect 14648 15076 14724 15110
rect 14539 15038 14724 15076
rect 14539 15004 14614 15038
rect 14648 15004 14724 15038
rect 14539 14966 14724 15004
rect 14539 14932 14614 14966
rect 14648 14932 14724 14966
rect 14029 14908 14170 14932
rect 245 14863 320 14897
rect 354 14863 430 14897
tri 792 14894 806 14908 ne
rect 806 14894 14170 14908
tri 14170 14894 14208 14932 nw
rect 14539 14894 14724 14932
rect 245 14825 430 14863
tri 806 14860 840 14894 ne
rect 840 14860 14136 14894
tri 14136 14860 14170 14894 nw
rect 14539 14860 14614 14894
rect 14648 14860 14724 14894
tri 840 14843 857 14860 ne
rect 857 14843 14119 14860
tri 14119 14843 14136 14860 nw
rect 245 14791 320 14825
rect 354 14791 430 14825
rect 245 14753 430 14791
rect 245 14719 320 14753
rect 354 14719 430 14753
rect 245 14681 430 14719
rect 245 14647 320 14681
rect 354 14647 430 14681
rect 245 14528 430 14647
rect 858 14774 2096 14843
rect 858 14740 883 14774
rect 917 14740 955 14774
rect 989 14740 1027 14774
rect 1061 14740 1099 14774
rect 1133 14740 1171 14774
rect 1205 14740 1243 14774
rect 1277 14740 1315 14774
rect 1349 14740 1387 14774
rect 1421 14740 1459 14774
rect 1493 14740 1531 14774
rect 1565 14740 1603 14774
rect 1637 14740 1675 14774
rect 1709 14740 1747 14774
rect 1781 14740 1819 14774
rect 1853 14740 1891 14774
rect 1925 14740 1963 14774
rect 1997 14740 2035 14774
rect 2069 14740 2096 14774
rect 858 14731 2096 14740
rect 245 14452 720 14528
rect 245 14418 320 14452
rect 354 14418 610 14452
rect 644 14418 720 14452
rect 245 14343 720 14418
rect 858 14295 908 14731
rect 2048 14295 2096 14731
rect 12858 14774 14096 14843
rect 12858 14740 12883 14774
rect 12917 14740 12955 14774
rect 12989 14740 13027 14774
rect 13061 14740 13099 14774
rect 13133 14740 13171 14774
rect 13205 14740 13243 14774
rect 13277 14740 13315 14774
rect 13349 14740 13387 14774
rect 13421 14740 13459 14774
rect 13493 14740 13531 14774
rect 13565 14740 13603 14774
rect 13637 14740 13675 14774
rect 13709 14740 13747 14774
rect 13781 14740 13819 14774
rect 13853 14740 13891 14774
rect 13925 14740 13963 14774
rect 13997 14740 14035 14774
rect 14069 14740 14096 14774
rect 12858 14731 14096 14740
rect 2248 14452 12705 14528
rect 2248 14418 2311 14452
rect 2345 14418 2383 14452
rect 2417 14418 2455 14452
rect 2489 14418 2527 14452
rect 2561 14418 2599 14452
rect 2633 14418 2671 14452
rect 2705 14418 2743 14452
rect 2777 14418 2815 14452
rect 2849 14418 2887 14452
rect 2921 14418 2959 14452
rect 2993 14418 3031 14452
rect 3065 14418 3103 14452
rect 3137 14418 3175 14452
rect 3209 14418 3247 14452
rect 3281 14418 3319 14452
rect 3353 14418 3391 14452
rect 3425 14418 3463 14452
rect 3497 14418 3535 14452
rect 3569 14418 3607 14452
rect 3641 14418 3679 14452
rect 3713 14418 3751 14452
rect 3785 14418 3823 14452
rect 3857 14418 3895 14452
rect 3929 14418 3967 14452
rect 4001 14418 4039 14452
rect 4073 14418 4111 14452
rect 4145 14418 4183 14452
rect 4217 14418 4255 14452
rect 4289 14418 4327 14452
rect 4361 14418 4399 14452
rect 4433 14418 4471 14452
rect 4505 14418 4543 14452
rect 4577 14418 4615 14452
rect 4649 14418 4687 14452
rect 4721 14418 4759 14452
rect 4793 14418 4831 14452
rect 4865 14418 4903 14452
rect 4937 14418 4975 14452
rect 5009 14418 5047 14452
rect 5081 14418 5119 14452
rect 5153 14418 5191 14452
rect 5225 14418 5263 14452
rect 5297 14418 5335 14452
rect 5369 14418 5407 14452
rect 5441 14418 5479 14452
rect 5513 14418 5551 14452
rect 5585 14418 5623 14452
rect 5657 14418 5695 14452
rect 5729 14418 5767 14452
rect 5801 14418 5839 14452
rect 5873 14418 5911 14452
rect 5945 14418 5983 14452
rect 6017 14418 6055 14452
rect 6089 14418 6127 14452
rect 6161 14418 6199 14452
rect 6233 14418 6271 14452
rect 6305 14418 6343 14452
rect 6377 14418 6415 14452
rect 6449 14418 6487 14452
rect 6521 14418 6559 14452
rect 6593 14418 6631 14452
rect 6665 14418 6703 14452
rect 6737 14418 6775 14452
rect 6809 14418 6847 14452
rect 6881 14418 6919 14452
rect 6953 14418 6991 14452
rect 7025 14418 7063 14452
rect 7097 14418 7135 14452
rect 7169 14418 7207 14452
rect 7241 14418 7279 14452
rect 7313 14418 7351 14452
rect 7385 14418 7423 14452
rect 7457 14418 7495 14452
rect 7529 14418 7567 14452
rect 7601 14418 7639 14452
rect 7673 14418 7711 14452
rect 7745 14418 7783 14452
rect 7817 14418 7855 14452
rect 7889 14418 7927 14452
rect 7961 14418 7999 14452
rect 8033 14418 8071 14452
rect 8105 14418 8143 14452
rect 8177 14418 8215 14452
rect 8249 14418 8287 14452
rect 8321 14418 8359 14452
rect 8393 14418 8431 14452
rect 8465 14418 8503 14452
rect 8537 14418 8575 14452
rect 8609 14418 8647 14452
rect 8681 14418 8719 14452
rect 8753 14418 8791 14452
rect 8825 14418 8863 14452
rect 8897 14418 8935 14452
rect 8969 14418 9007 14452
rect 9041 14418 9079 14452
rect 9113 14418 9151 14452
rect 9185 14418 9223 14452
rect 9257 14418 9295 14452
rect 9329 14418 9367 14452
rect 9401 14418 9439 14452
rect 9473 14418 9511 14452
rect 9545 14418 9583 14452
rect 9617 14418 9655 14452
rect 9689 14418 9727 14452
rect 9761 14418 9799 14452
rect 9833 14418 9871 14452
rect 9905 14418 9943 14452
rect 9977 14418 10015 14452
rect 10049 14418 10087 14452
rect 10121 14418 10159 14452
rect 10193 14418 10231 14452
rect 10265 14418 10303 14452
rect 10337 14418 10375 14452
rect 10409 14418 10447 14452
rect 10481 14418 10519 14452
rect 10553 14418 10591 14452
rect 10625 14418 10663 14452
rect 10697 14418 10735 14452
rect 10769 14418 10807 14452
rect 10841 14418 10879 14452
rect 10913 14418 10951 14452
rect 10985 14418 11023 14452
rect 11057 14418 11095 14452
rect 11129 14418 11167 14452
rect 11201 14418 11239 14452
rect 11273 14418 11311 14452
rect 11345 14418 11383 14452
rect 11417 14418 11455 14452
rect 11489 14418 11527 14452
rect 11561 14418 11599 14452
rect 11633 14418 11671 14452
rect 11705 14418 11743 14452
rect 11777 14418 11815 14452
rect 11849 14418 11887 14452
rect 11921 14418 11959 14452
rect 11993 14418 12031 14452
rect 12065 14418 12103 14452
rect 12137 14418 12175 14452
rect 12209 14418 12247 14452
rect 12281 14418 12319 14452
rect 12353 14418 12391 14452
rect 12425 14418 12463 14452
rect 12497 14418 12535 14452
rect 12569 14418 12607 14452
rect 12641 14418 12705 14452
rect 2248 14343 12705 14418
rect 858 14252 2096 14295
rect 12858 14295 12908 14731
rect 14048 14295 14096 14731
rect 14539 14822 14724 14860
rect 14539 14788 14614 14822
rect 14648 14788 14724 14822
rect 14539 14750 14724 14788
rect 14539 14716 14614 14750
rect 14648 14716 14724 14750
rect 14539 14678 14724 14716
rect 14539 14644 14614 14678
rect 14648 14644 14724 14678
rect 14539 14528 14724 14644
rect 14232 14452 14724 14528
rect 14232 14418 14314 14452
rect 14348 14418 14614 14452
rect 14648 14418 14724 14452
rect 14232 14343 14724 14418
rect 12858 14252 14096 14295
<< via1 >>
rect 957 36498 2161 37211
rect 12821 36498 14025 37208
rect 957 36464 988 36498
rect 988 36464 1022 36498
rect 1022 36464 1060 36498
rect 1060 36464 1094 36498
rect 1094 36464 1132 36498
rect 1132 36464 1166 36498
rect 1166 36464 1204 36498
rect 1204 36464 1238 36498
rect 1238 36464 1276 36498
rect 1276 36464 1310 36498
rect 1310 36464 1348 36498
rect 1348 36464 1382 36498
rect 1382 36464 1420 36498
rect 1420 36464 1454 36498
rect 1454 36464 1492 36498
rect 1492 36464 1526 36498
rect 1526 36464 1564 36498
rect 1564 36464 1598 36498
rect 1598 36464 1636 36498
rect 1636 36464 1670 36498
rect 1670 36464 1708 36498
rect 1708 36464 1742 36498
rect 1742 36464 1780 36498
rect 1780 36464 1814 36498
rect 1814 36464 1852 36498
rect 1852 36464 1886 36498
rect 1886 36464 1924 36498
rect 1924 36464 1958 36498
rect 1958 36464 1996 36498
rect 1996 36464 2030 36498
rect 2030 36464 2068 36498
rect 2068 36464 2102 36498
rect 2102 36464 2140 36498
rect 2140 36464 2161 36498
rect 12821 36464 12830 36498
rect 12830 36464 12868 36498
rect 12868 36464 12902 36498
rect 12902 36464 12940 36498
rect 12940 36464 12974 36498
rect 12974 36464 13012 36498
rect 13012 36464 13046 36498
rect 13046 36464 13084 36498
rect 13084 36464 13118 36498
rect 13118 36464 13156 36498
rect 13156 36464 13190 36498
rect 13190 36464 13228 36498
rect 13228 36464 13262 36498
rect 13262 36464 13300 36498
rect 13300 36464 13334 36498
rect 13334 36464 13372 36498
rect 13372 36464 13406 36498
rect 13406 36464 13444 36498
rect 13444 36464 13478 36498
rect 13478 36464 13516 36498
rect 13516 36464 13550 36498
rect 13550 36464 13588 36498
rect 13588 36464 13622 36498
rect 13622 36464 13660 36498
rect 13660 36464 13694 36498
rect 13694 36464 13732 36498
rect 13732 36464 13766 36498
rect 13766 36464 13804 36498
rect 13804 36464 13838 36498
rect 13838 36464 13876 36498
rect 13876 36464 13910 36498
rect 13910 36464 13948 36498
rect 13948 36464 13982 36498
rect 13982 36464 14020 36498
rect 14020 36464 14025 36498
rect 957 36455 2161 36464
rect 12821 36452 14025 36464
rect 4944 29407 7236 30227
rect 7745 29407 10037 30227
rect 4939 28219 7231 28335
rect 7750 28219 10042 28335
rect 2509 27906 4481 28022
rect 10500 27906 12472 28022
rect 4939 27603 7231 27719
rect 7750 27603 10042 27719
rect 4933 25909 7225 26025
rect 7757 25909 10049 26025
rect 2546 25643 4454 25759
rect 10528 25643 12436 25759
rect 4933 25377 7225 25493
rect 7757 25377 10049 25493
rect 4945 23669 7237 24489
rect 7744 23669 10036 24489
rect 908 14295 2048 14731
rect 12908 14295 14048 14731
<< metal2 >>
tri 4891 39322 4991 39422 se
rect 4991 39322 7191 39422
tri 7191 39322 7291 39422 sw
rect 4891 39213 7291 39322
rect 885 37211 2234 37258
rect 885 36455 957 37211
rect 2161 36455 2234 37211
rect 885 36408 2234 36455
rect 4891 35317 4979 39213
rect 7195 35317 7291 39213
rect 4891 30227 7291 35317
rect 4891 29407 4944 30227
rect 7236 29407 7291 30227
tri 301 28975 501 29175 se
rect 501 28975 4291 29175
tri 4291 28975 4491 29175 sw
rect 301 28859 4491 28975
rect 301 24803 466 28859
rect 2442 28022 4491 28859
rect 2442 27906 2509 28022
rect 4481 27906 4491 28022
rect 2442 25759 4491 27906
rect 4891 28335 7291 29407
rect 4891 28219 4939 28335
rect 7231 28219 7291 28335
rect 4891 27719 7291 28219
rect 4891 27603 4939 27719
rect 7231 27603 7291 27719
rect 4891 27317 7291 27603
tri 4891 27117 5091 27317 ne
rect 5091 27117 7091 27317
tri 7091 27117 7291 27317 nw
tri 7691 39322 7791 39422 se
rect 7791 39322 9991 39422
tri 9991 39322 10091 39422 sw
rect 7691 39213 10091 39322
rect 7691 35317 7779 39213
rect 9995 35317 10091 39213
rect 12752 37208 14101 37262
rect 12752 36452 12821 37208
rect 14025 36452 14101 37208
rect 12752 36412 14101 36452
rect 7691 30227 10091 35317
rect 7691 29407 7745 30227
rect 10037 29407 10091 30227
rect 7691 28335 10091 29407
rect 7691 28219 7750 28335
rect 10042 28219 10091 28335
rect 7691 27719 10091 28219
rect 7691 27603 7750 27719
rect 10042 27603 10091 27719
rect 7691 27317 10091 27603
tri 7691 27117 7891 27317 ne
rect 7891 27117 9891 27317
tri 9891 27117 10091 27317 nw
tri 10491 28975 10691 29175 se
rect 10691 28975 14431 29175
tri 14431 28975 14631 29175 sw
rect 10491 28907 14631 28975
rect 10491 28022 12455 28907
rect 10491 27906 10500 28022
rect 2442 25643 2546 25759
rect 4454 25643 4491 25759
rect 2442 24803 4491 25643
rect 301 24516 4491 24803
tri 301 24503 314 24516 ne
rect 314 24503 4478 24516
tri 4478 24503 4491 24516 nw
tri 4891 26278 5091 26478 se
rect 5091 26278 7091 26478
tri 7091 26278 7291 26478 sw
rect 4891 26025 7291 26278
rect 4891 25909 4933 26025
rect 7225 25909 7291 26025
rect 4891 25493 7291 25909
rect 4891 25377 4933 25493
rect 7225 25377 7291 25493
tri 314 24489 328 24503 ne
rect 328 24489 4464 24503
tri 4464 24489 4478 24503 nw
rect 4891 24489 7291 25377
tri 328 24316 501 24489 ne
rect 501 24316 4291 24489
tri 4291 24316 4464 24489 nw
rect 4891 23669 4945 24489
rect 7237 23669 7291 24489
tri 2891 19364 4891 21364 se
rect 4891 19364 7291 23669
rect 2891 18931 5291 19364
rect 2891 17275 2942 18931
rect 5238 17275 5291 18931
tri 5291 17364 7291 19364 nw
tri 7691 26278 7891 26478 se
rect 7891 26278 9891 26478
tri 9891 26278 10091 26478 sw
rect 7691 26025 10091 26278
rect 7691 25909 7757 26025
rect 10049 25909 10091 26025
rect 7691 25493 10091 25909
rect 7691 25377 7757 25493
rect 10049 25377 10091 25493
rect 7691 24489 10091 25377
rect 7691 23669 7744 24489
rect 10036 23669 10091 24489
rect 10491 25759 12455 27906
rect 10491 25643 10528 25759
rect 12436 25643 12455 25759
rect 10491 24851 12455 25643
rect 14431 24851 14631 28907
rect 10491 24516 14631 24851
tri 10491 24316 10691 24516 ne
rect 10691 24316 14431 24516
tri 14431 24316 14631 24516 nw
rect 7691 19330 10091 23669
tri 10091 19330 12091 21330 sw
tri 7691 17364 9657 19330 ne
rect 9657 18931 12091 19330
rect 9657 17364 9742 18931
tri 9657 17330 9691 17364 ne
rect 2891 17214 5291 17275
rect 2891 17086 3103 17214
tri 2891 16986 2991 17086 ne
rect 2991 17078 3103 17086
rect 5239 17078 5291 17214
rect 2991 17056 5291 17078
rect 2991 16986 5221 17056
tri 5221 16986 5291 17056 nw
rect 9691 17275 9742 17364
rect 12038 17275 12091 18931
rect 9691 17214 12091 17275
rect 9691 17078 9739 17214
rect 11875 17086 12091 17214
rect 11875 17078 11991 17086
rect 9691 17056 11991 17078
tri 9691 16986 9761 17056 ne
rect 9761 16986 11991 17056
tri 11991 16986 12091 17086 nw
rect 858 14731 2096 14772
rect 858 14295 908 14731
rect 2048 14295 2096 14731
rect 858 14252 2096 14295
rect 12858 14731 14096 14772
rect 12858 14295 12908 14731
rect 14048 14295 14096 14731
rect 12858 14252 14096 14295
<< via2 >>
rect 971 36485 2147 37181
rect 4979 35317 7195 39213
rect 466 24803 2442 28859
rect 7779 35317 9995 39213
rect 12835 36482 14011 37178
rect 12455 28022 14431 28907
rect 12455 27906 12472 28022
rect 12472 27906 14431 28022
rect 2942 17275 5238 18931
rect 12455 24851 14431 27906
rect 3103 17078 5239 17214
rect 9742 17275 12038 18931
rect 9739 17078 11875 17214
<< metal3 >>
tri 4805 39522 5205 39922 se
rect 5205 39857 9786 39922
rect 5205 39553 5267 39857
rect 9731 39553 9786 39857
rect 5205 39522 9786 39553
tri 9786 39522 10186 39922 sw
rect 4805 39455 10186 39522
rect 885 37185 2234 37258
rect 885 36481 967 37185
rect 2151 36481 2234 37185
rect 885 36408 2234 36481
rect 4805 35311 4975 39455
rect 9999 35311 10186 39455
rect 12752 37182 14101 37262
rect 12752 36478 12831 37182
rect 14015 36478 14101 37182
rect 12752 36412 14101 36478
rect 4805 35266 10186 35311
tri 4805 35166 4905 35266 ne
rect 4905 35166 10086 35266
tri 10086 35166 10186 35266 nw
tri 245 33721 1155 34631 se
rect 1155 34575 3100 34631
rect 1155 34111 2339 34575
rect 3043 34111 3100 34575
rect 1155 33848 3100 34111
rect 1155 33721 2700 33848
rect 245 32961 2700 33721
tri 2700 33448 3100 33848 nw
rect 11900 34574 13835 34631
rect 11900 34110 11969 34574
rect 12673 34110 13835 34574
rect 11900 33848 13835 34110
tri 11900 33448 12300 33848 ne
rect 12300 33742 13835 33848
tri 13835 33742 14724 34631 sw
rect 245 28859 1043 32961
rect 1427 28859 2700 32961
rect 245 24803 466 28859
rect 2442 24803 2700 28859
rect 245 21217 1043 24803
rect 1427 21217 2700 24803
rect 245 20438 2700 21217
tri 245 19528 1155 20438 ne
rect 1155 20067 2700 20438
rect 12300 32853 14724 33742
rect 12300 28907 13589 32853
rect 13973 28907 14724 32853
rect 12300 24851 12455 28907
rect 14431 24851 14724 28907
rect 12300 21109 13589 24851
rect 13973 21109 14724 24851
rect 12300 20448 14724 21109
tri 2700 20067 2912 20279 sw
tri 12108 20067 12300 20259 se
rect 12300 20067 13804 20448
rect 1155 20027 13804 20067
rect 1155 19563 2316 20027
rect 12700 19563 13804 20027
rect 1155 19528 13804 19563
tri 13804 19528 14724 20448 nw
tri 2842 18996 3042 19196 se
rect 3042 18996 5380 19196
rect 2842 18931 5380 18996
rect 2842 18895 2942 18931
rect 5238 18895 5380 18931
rect 2842 17311 2938 18895
rect 5242 17311 5380 18895
rect 2842 17275 2942 17311
rect 5238 17275 5380 17311
rect 2842 17230 5380 17275
tri 2842 17214 2858 17230 ne
rect 2858 17218 5380 17230
rect 2858 17214 3099 17218
tri 2858 17078 2994 17214 ne
rect 2994 17078 3099 17214
tri 2994 17061 3011 17078 ne
rect 3011 17074 3099 17078
rect 5243 17074 5380 17218
rect 3011 17061 5380 17074
tri 3011 17030 3042 17061 ne
rect 3042 17030 5380 17061
rect 9596 18996 11935 19196
tri 11935 18996 12135 19196 sw
rect 9596 18931 12135 18996
rect 9596 18895 9742 18931
rect 12038 18895 12135 18931
rect 9596 17311 9738 18895
rect 12042 17311 12135 18895
rect 9596 17275 9742 17311
rect 12038 17275 12135 17311
rect 9596 17230 12135 17275
rect 9596 17218 11935 17230
rect 9596 17074 9735 17218
rect 11879 17074 11935 17218
rect 9596 17030 11935 17074
tri 11935 17030 12135 17230 nw
rect 858 14705 2096 14772
rect 858 14321 926 14705
rect 2030 14321 2096 14705
rect 858 14252 2096 14321
rect 12858 14705 14096 14772
rect 12858 14321 12926 14705
rect 14030 14321 14096 14705
rect 12858 14252 14096 14321
<< via3 >>
rect 5267 39553 9731 39857
rect 967 37181 2151 37185
rect 967 36485 971 37181
rect 971 36485 2147 37181
rect 2147 36485 2151 37181
rect 967 36481 2151 36485
rect 4975 39213 9999 39455
rect 4975 35317 4979 39213
rect 4979 35317 7195 39213
rect 7195 35317 7779 39213
rect 7779 35317 9995 39213
rect 9995 35317 9999 39213
rect 4975 35311 9999 35317
rect 12831 37178 14015 37182
rect 12831 36482 12835 37178
rect 12835 36482 14011 37178
rect 14011 36482 14015 37178
rect 12831 36478 14015 36482
rect 2339 34111 3043 34575
rect 11969 34110 12673 34574
rect 1043 28859 1427 32961
rect 1043 24803 1427 28859
rect 1043 21217 1427 24803
rect 13589 28907 13973 32853
rect 13589 24851 13973 28907
rect 13589 21109 13973 24851
rect 2316 19563 12700 20027
rect 2938 17311 2942 18895
rect 2942 17311 5238 18895
rect 5238 17311 5242 18895
rect 3099 17214 5243 17218
rect 3099 17078 3103 17214
rect 3103 17078 5239 17214
rect 5239 17078 5243 17214
rect 3099 17074 5243 17078
rect 9738 17311 9742 18895
rect 9742 17311 12038 18895
rect 12038 17311 12042 18895
rect 9735 17214 11879 17218
rect 9735 17078 9739 17214
rect 9739 17078 11875 17214
rect 11875 17078 11879 17214
rect 9735 17074 11879 17078
rect 926 14321 2030 14705
rect 12926 14321 14030 14705
<< metal4 >>
rect 8 35144 262 39987
rect 5257 39857 9742 39861
rect 5257 39553 5267 39857
rect 9731 39553 9742 39857
rect 5257 39550 9742 39553
rect 4949 39455 10025 39476
rect 932 37185 2187 37214
rect 932 36481 967 37185
rect 2151 36481 2187 37185
rect 932 36453 2187 36481
rect 4949 35311 4975 39455
rect 9999 35311 10025 39455
rect 12796 37182 14051 37211
rect 12796 36478 12831 37182
rect 14015 36478 14051 37182
rect 12796 36450 14051 36478
rect 4949 35290 10025 35311
rect 14754 35144 15008 39987
rect 2305 34575 3078 34591
rect 2305 34111 2339 34575
rect 3043 34111 3078 34575
rect 2305 34096 3078 34111
rect 11935 34574 12708 34590
rect 11935 34110 11969 34574
rect 12673 34110 12708 34574
rect 11935 34095 12708 34110
rect 1004 32961 1466 32980
rect 1004 21217 1043 32961
rect 1427 21217 1466 32961
rect 1004 21198 1466 21217
rect 13550 32853 14012 32872
rect 13550 21109 13589 32853
rect 13973 21109 14012 32853
rect 13550 21090 14012 21109
rect 2299 20027 12718 20035
rect 2299 19563 2316 20027
rect 12700 19563 12718 20027
rect 2299 19555 12718 19563
tri 6512 19127 6912 19527 ne
rect 8 13994 262 18987
rect 2912 18895 5268 18934
rect 2912 17311 2938 18895
rect 5242 17311 5268 18895
rect 2912 17273 5268 17311
rect 3077 17218 5265 17231
rect 3077 17074 3099 17218
rect 5243 17074 5265 17218
rect 3077 17061 5265 17074
rect 908 14705 2048 14731
rect 908 14321 926 14705
rect 2030 14321 2048 14705
rect 908 14295 2048 14321
rect 6912 13996 8112 19528
tri 8112 19127 8512 19527 nw
rect 9712 18895 12068 18934
rect 9712 17311 9738 18895
rect 12042 17311 12068 18895
rect 9712 17273 12068 17311
rect 9713 17218 11901 17231
rect 9713 17074 9735 17218
rect 11879 17074 11901 17218
rect 9713 17061 11901 17074
rect 12908 14705 14048 14731
rect 12908 14321 12926 14705
rect 14030 14321 14048 14705
rect 12908 14295 14048 14321
rect 14754 13994 15008 18987
use sky130_ef_io__com_pg_esd  sky130_ef_io__com_pg_esd_0
timestamp 1686671242
transform 1 0 0 0 1 0
box 8 13994 15008 39987
use sky130_ef_io__esd_ndiode_11v0_single  sky130_ef_io__minesd_vddio
timestamp 1686671242
transform 0 1 7496 -1 0 26758
box 160 -5766 1962 5766
use sky130_ef_io__esd_pdiode_11v0_single  sky130_ef_io__minesd_vssio
timestamp 1686671242
transform 0 1 7508 -1 0 29198
box 896 -5188 1566 5188
<< labels >>
flabel metal4 s 14754 35144 15008 39987 3 FreeSans 650 180 0 0 sky130_fd_io__com_bus_hookup_0.VSSIO
flabel metal4 s 14754 13994 15008 18987 3 FreeSans 650 180 0 0 sky130_fd_io__com_bus_hookup_0.VDDIO
flabel metal4 s 8 35144 262 39987 3 FreeSans 650 0 0 0 sky130_fd_io__com_bus_hookup_0.VSSIO
flabel metal4 s 8 13994 262 18987 3 FreeSans 650 0 0 0 sky130_fd_io__com_bus_hookup_0.VDDIO
flabel metal4 s 6912 13996 8112 14196 0 FreeSans 1400 0 0 0 P_CORE
port 1 nsew
<< properties >>
string GDS_END 7522862
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 5766234
<< end >>
