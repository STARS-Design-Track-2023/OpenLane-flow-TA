magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 3 21 549 203
rect 29 -17 63 21
<< scnmos >>
rect 81 47 111 177
rect 269 47 299 177
rect 354 47 384 177
rect 440 47 470 177
<< scpmoshvt >>
rect 81 297 111 497
rect 269 297 299 497
rect 354 297 384 497
rect 440 297 470 497
<< ndiff >>
rect 29 129 81 177
rect 29 95 37 129
rect 71 95 81 129
rect 29 47 81 95
rect 111 89 269 177
rect 111 55 139 89
rect 173 55 207 89
rect 241 55 269 89
rect 111 47 269 55
rect 299 127 354 177
rect 299 93 309 127
rect 343 93 354 127
rect 299 47 354 93
rect 384 47 440 177
rect 470 123 523 177
rect 470 89 481 123
rect 515 89 523 123
rect 470 47 523 89
<< pdiff >>
rect 29 459 81 497
rect 29 425 37 459
rect 71 425 81 459
rect 29 371 81 425
rect 29 337 37 371
rect 71 337 81 371
rect 29 297 81 337
rect 111 485 163 497
rect 111 451 121 485
rect 155 451 163 485
rect 111 417 163 451
rect 111 383 121 417
rect 155 383 163 417
rect 111 297 163 383
rect 217 453 269 497
rect 217 419 225 453
rect 259 419 269 453
rect 217 379 269 419
rect 217 345 225 379
rect 259 345 269 379
rect 217 297 269 345
rect 299 457 354 497
rect 299 423 309 457
rect 343 423 354 457
rect 299 383 354 423
rect 299 349 309 383
rect 343 349 354 383
rect 299 297 354 349
rect 384 489 440 497
rect 384 455 395 489
rect 429 455 440 489
rect 384 421 440 455
rect 384 387 395 421
rect 429 387 440 421
rect 384 297 440 387
rect 470 457 523 497
rect 470 423 481 457
rect 515 423 523 457
rect 470 383 523 423
rect 470 349 481 383
rect 515 349 523 383
rect 470 297 523 349
<< ndiffc >>
rect 37 95 71 129
rect 139 55 173 89
rect 207 55 241 89
rect 309 93 343 127
rect 481 89 515 123
<< pdiffc >>
rect 37 425 71 459
rect 37 337 71 371
rect 121 451 155 485
rect 121 383 155 417
rect 225 419 259 453
rect 225 345 259 379
rect 309 423 343 457
rect 309 349 343 383
rect 395 455 429 489
rect 395 387 429 421
rect 481 423 515 457
rect 481 349 515 383
<< poly >>
rect 81 497 111 523
rect 269 497 299 523
rect 354 497 384 523
rect 440 497 470 523
rect 81 265 111 297
rect 269 265 299 297
rect 354 265 384 297
rect 440 265 470 297
rect 81 249 166 265
rect 81 215 122 249
rect 156 215 166 249
rect 81 199 166 215
rect 214 249 299 265
rect 214 215 224 249
rect 258 215 299 249
rect 214 199 299 215
rect 342 249 396 265
rect 342 215 352 249
rect 386 215 396 249
rect 342 199 396 215
rect 440 249 524 265
rect 440 215 480 249
rect 514 215 524 249
rect 440 199 524 215
rect 81 177 111 199
rect 269 177 299 199
rect 354 177 384 199
rect 440 177 470 199
rect 81 21 111 47
rect 269 21 299 47
rect 354 21 384 47
rect 440 21 470 47
<< polycont >>
rect 122 215 156 249
rect 224 215 258 249
rect 352 215 386 249
rect 480 215 514 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 19 459 71 491
rect 19 425 37 459
rect 19 371 71 425
rect 105 485 173 527
rect 105 451 121 485
rect 155 451 173 485
rect 105 417 173 451
rect 105 383 121 417
rect 155 383 173 417
rect 105 381 173 383
rect 209 453 263 491
rect 209 419 225 453
rect 259 419 263 453
rect 19 337 37 371
rect 209 379 263 419
rect 209 345 225 379
rect 259 345 263 379
rect 19 129 71 337
rect 19 95 37 129
rect 109 301 263 345
rect 299 457 345 491
rect 299 423 309 457
rect 343 423 345 457
rect 299 383 345 423
rect 379 489 445 527
rect 379 455 395 489
rect 429 455 445 489
rect 379 421 445 455
rect 379 387 395 421
rect 429 387 445 421
rect 379 385 445 387
rect 479 457 531 491
rect 479 423 481 457
rect 515 423 531 457
rect 299 349 309 383
rect 343 349 345 383
rect 479 383 531 423
rect 479 349 481 383
rect 515 349 531 383
rect 299 301 531 349
rect 109 249 167 301
rect 109 215 122 249
rect 156 215 167 249
rect 109 167 167 215
rect 203 249 296 265
rect 203 215 224 249
rect 258 215 296 249
rect 203 203 296 215
rect 332 249 437 265
rect 332 215 352 249
rect 386 215 437 249
rect 332 203 437 215
rect 109 127 355 167
rect 19 53 71 95
rect 293 93 309 127
rect 343 93 355 127
rect 123 89 257 91
rect 123 55 139 89
rect 173 55 207 89
rect 241 55 257 89
rect 123 17 257 55
rect 293 53 355 93
rect 391 75 437 203
rect 473 249 533 265
rect 473 215 480 249
rect 514 215 533 249
rect 473 199 533 215
rect 473 123 531 163
rect 473 89 481 123
rect 515 89 531 123
rect 473 17 531 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 397 85 431 119 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 397 153 431 187 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 29 85 63 119 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 29 425 63 459 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 29 357 63 391 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a21o_1
rlabel metal1 s 0 -48 552 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 4032030
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4026040
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 13.800 13.600 
<< end >>
