magic
tech sky130A
magscale 1 2
timestamp 1686671242
<< pwell >>
rect 15 163 787 817
<< nmoslvt >>
rect 171 189 201 791
rect 257 189 287 791
rect 343 189 373 791
rect 429 189 459 791
rect 515 189 545 791
rect 601 189 631 791
<< ndiff >>
rect 111 779 171 791
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 779 257 791
rect 201 513 212 779
rect 246 513 257 779
rect 201 467 257 513
rect 201 201 212 467
rect 246 201 257 467
rect 201 189 257 201
rect 287 779 343 791
rect 287 513 298 779
rect 332 513 343 779
rect 287 467 343 513
rect 287 201 298 467
rect 332 201 343 467
rect 287 189 343 201
rect 373 779 429 791
rect 373 513 384 779
rect 418 513 429 779
rect 373 467 429 513
rect 373 201 384 467
rect 418 201 429 467
rect 373 189 429 201
rect 459 779 515 791
rect 459 513 470 779
rect 504 513 515 779
rect 459 467 515 513
rect 459 201 470 467
rect 504 201 515 467
rect 459 189 515 201
rect 545 779 601 791
rect 545 513 556 779
rect 590 513 601 779
rect 545 467 601 513
rect 545 201 556 467
rect 590 201 601 467
rect 545 189 601 201
rect 631 779 691 791
rect 631 745 642 779
rect 676 745 691 779
rect 631 711 691 745
rect 631 677 642 711
rect 676 677 691 711
rect 631 643 691 677
rect 631 609 642 643
rect 676 609 691 643
rect 631 575 691 609
rect 631 541 642 575
rect 676 541 691 575
rect 631 507 691 541
rect 631 473 642 507
rect 676 473 691 507
rect 631 439 691 473
rect 631 405 642 439
rect 676 405 691 439
rect 631 371 691 405
rect 631 337 642 371
rect 676 337 691 371
rect 631 303 691 337
rect 631 269 642 303
rect 676 269 691 303
rect 631 235 691 269
rect 631 201 642 235
rect 676 201 691 235
rect 631 189 691 201
<< ndiffc >>
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 513 246 779
rect 212 201 246 467
rect 298 513 332 779
rect 298 201 332 467
rect 384 513 418 779
rect 384 201 418 467
rect 470 513 504 779
rect 470 201 504 467
rect 556 513 590 779
rect 556 201 590 467
rect 642 745 676 779
rect 642 677 676 711
rect 642 609 676 643
rect 642 541 676 575
rect 642 473 676 507
rect 642 405 676 439
rect 642 337 676 371
rect 642 269 676 303
rect 642 201 676 235
<< psubdiff >>
rect 41 779 111 791
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 691 779 761 791
rect 691 745 710 779
rect 744 745 761 779
rect 691 711 761 745
rect 691 677 710 711
rect 744 677 761 711
rect 691 643 761 677
rect 691 609 710 643
rect 744 609 761 643
rect 691 575 761 609
rect 691 541 710 575
rect 744 541 761 575
rect 691 507 761 541
rect 691 473 710 507
rect 744 473 761 507
rect 691 439 761 473
rect 691 405 710 439
rect 744 405 761 439
rect 691 371 761 405
rect 691 337 710 371
rect 744 337 761 371
rect 691 303 761 337
rect 691 269 710 303
rect 744 269 761 303
rect 691 235 761 269
rect 691 201 710 235
rect 744 201 761 235
rect 691 189 761 201
<< psubdiffcont >>
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 710 745 744 779
rect 710 677 744 711
rect 710 609 744 643
rect 710 541 744 575
rect 710 473 744 507
rect 710 405 744 439
rect 710 337 744 371
rect 710 269 744 303
rect 710 201 744 235
<< poly >>
rect 243 891 559 907
rect 120 867 201 883
rect 120 833 136 867
rect 170 833 201 867
rect 243 857 264 891
rect 538 857 559 891
rect 243 841 559 857
rect 601 867 682 883
rect 120 817 201 833
rect 171 791 201 817
rect 257 791 287 841
rect 343 791 373 841
rect 429 791 459 841
rect 515 791 545 841
rect 601 833 632 867
rect 666 833 682 867
rect 601 817 682 833
rect 601 791 631 817
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 287 189
rect 343 139 373 189
rect 429 139 459 189
rect 515 139 545 189
rect 601 163 631 189
rect 601 147 682 163
rect 120 97 201 113
rect 243 123 559 139
rect 243 89 264 123
rect 538 89 559 123
rect 601 113 632 147
rect 666 113 682 147
rect 601 97 682 113
rect 243 73 559 89
<< polycont >>
rect 136 833 170 867
rect 264 857 538 891
rect 632 833 666 867
rect 136 113 170 147
rect 264 89 538 123
rect 632 113 666 147
<< locali >>
rect 243 961 559 980
rect 243 927 255 961
rect 289 927 337 961
rect 371 927 431 961
rect 465 927 513 961
rect 547 927 559 961
rect 243 891 559 927
rect 243 889 264 891
rect 538 889 559 891
rect 120 867 186 883
rect 120 833 136 867
rect 170 833 186 867
rect 243 855 255 889
rect 289 855 337 857
rect 371 855 431 857
rect 465 855 513 857
rect 547 855 559 889
rect 243 841 559 855
rect 616 867 682 883
rect 120 817 186 833
rect 616 833 632 867
rect 666 833 682 867
rect 616 817 682 833
rect 120 795 160 817
rect 642 795 682 817
rect 41 779 160 795
rect 41 745 58 779
rect 92 759 126 779
rect 94 745 126 759
rect 41 725 60 745
rect 94 725 160 745
rect 41 711 160 725
rect 41 677 58 711
rect 92 687 126 711
rect 94 677 126 687
rect 41 653 60 677
rect 94 653 160 677
rect 41 643 160 653
rect 41 609 58 643
rect 92 615 126 643
rect 94 609 126 615
rect 41 581 60 609
rect 94 581 160 609
rect 41 575 160 581
rect 41 541 58 575
rect 92 543 126 575
rect 94 541 126 543
rect 41 509 60 541
rect 94 509 160 541
rect 41 507 160 509
rect 41 473 58 507
rect 92 473 126 507
rect 41 471 160 473
rect 41 439 60 471
rect 94 439 160 471
rect 41 405 58 439
rect 94 437 126 439
rect 92 405 126 437
rect 41 399 160 405
rect 41 371 60 399
rect 94 371 160 399
rect 41 337 58 371
rect 94 365 126 371
rect 92 337 126 365
rect 41 327 160 337
rect 41 303 60 327
rect 94 303 160 327
rect 41 269 58 303
rect 94 293 126 303
rect 92 269 126 293
rect 41 255 160 269
rect 41 235 60 255
rect 94 235 160 255
rect 41 201 58 235
rect 94 221 126 235
rect 92 201 126 221
rect 41 185 160 201
rect 212 779 246 795
rect 212 471 246 509
rect 212 185 246 201
rect 298 779 332 795
rect 298 471 332 509
rect 298 185 332 201
rect 384 779 418 795
rect 384 471 418 509
rect 384 185 418 201
rect 470 779 504 795
rect 470 471 504 509
rect 470 185 504 201
rect 556 779 590 795
rect 556 471 590 509
rect 556 185 590 201
rect 642 779 761 795
rect 676 759 710 779
rect 676 745 708 759
rect 744 745 761 779
rect 642 725 708 745
rect 742 725 761 745
rect 642 711 761 725
rect 676 687 710 711
rect 676 677 708 687
rect 744 677 761 711
rect 642 653 708 677
rect 742 653 761 677
rect 642 643 761 653
rect 676 615 710 643
rect 676 609 708 615
rect 744 609 761 643
rect 642 581 708 609
rect 742 581 761 609
rect 642 575 761 581
rect 676 543 710 575
rect 676 541 708 543
rect 744 541 761 575
rect 642 509 708 541
rect 742 509 761 541
rect 642 507 761 509
rect 676 473 710 507
rect 744 473 761 507
rect 642 471 761 473
rect 642 439 708 471
rect 742 439 761 471
rect 676 437 708 439
rect 676 405 710 437
rect 744 405 761 439
rect 642 399 761 405
rect 642 371 708 399
rect 742 371 761 399
rect 676 365 708 371
rect 676 337 710 365
rect 744 337 761 371
rect 642 327 761 337
rect 642 303 708 327
rect 742 303 761 327
rect 676 293 708 303
rect 676 269 710 293
rect 744 269 761 303
rect 642 255 761 269
rect 642 235 708 255
rect 742 235 761 255
rect 676 221 708 235
rect 676 201 710 221
rect 744 201 761 235
rect 642 185 761 201
rect 120 163 160 185
rect 642 163 682 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 616 147 682 163
rect 120 97 186 113
rect 243 125 559 139
rect 243 91 255 125
rect 289 123 337 125
rect 371 123 431 125
rect 465 123 513 125
rect 547 91 559 125
rect 616 113 632 147
rect 666 113 682 147
rect 616 97 682 113
rect 243 89 264 91
rect 538 89 559 91
rect 243 53 559 89
rect 243 19 255 53
rect 289 19 337 53
rect 371 19 431 53
rect 465 19 513 53
rect 547 19 559 53
rect 243 0 559 19
<< viali >>
rect 255 927 289 961
rect 337 927 371 961
rect 431 927 465 961
rect 513 927 547 961
rect 255 857 264 889
rect 264 857 289 889
rect 337 857 371 889
rect 431 857 465 889
rect 513 857 538 889
rect 538 857 547 889
rect 255 855 289 857
rect 337 855 371 857
rect 431 855 465 857
rect 513 855 547 857
rect 60 745 92 759
rect 92 745 94 759
rect 60 725 94 745
rect 60 677 92 687
rect 92 677 94 687
rect 60 653 94 677
rect 60 609 92 615
rect 92 609 94 615
rect 60 581 94 609
rect 60 541 92 543
rect 92 541 94 543
rect 60 509 94 541
rect 60 439 94 471
rect 60 437 92 439
rect 92 437 94 439
rect 60 371 94 399
rect 60 365 92 371
rect 92 365 94 371
rect 60 303 94 327
rect 60 293 92 303
rect 92 293 94 303
rect 60 235 94 255
rect 60 221 92 235
rect 92 221 94 235
rect 212 725 246 759
rect 212 653 246 687
rect 212 581 246 615
rect 212 513 246 543
rect 212 509 246 513
rect 212 467 246 471
rect 212 437 246 467
rect 212 365 246 399
rect 212 293 246 327
rect 212 221 246 255
rect 298 725 332 759
rect 298 653 332 687
rect 298 581 332 615
rect 298 513 332 543
rect 298 509 332 513
rect 298 467 332 471
rect 298 437 332 467
rect 298 365 332 399
rect 298 293 332 327
rect 298 221 332 255
rect 384 725 418 759
rect 384 653 418 687
rect 384 581 418 615
rect 384 513 418 543
rect 384 509 418 513
rect 384 467 418 471
rect 384 437 418 467
rect 384 365 418 399
rect 384 293 418 327
rect 384 221 418 255
rect 470 725 504 759
rect 470 653 504 687
rect 470 581 504 615
rect 470 513 504 543
rect 470 509 504 513
rect 470 467 504 471
rect 470 437 504 467
rect 470 365 504 399
rect 470 293 504 327
rect 470 221 504 255
rect 556 725 590 759
rect 556 653 590 687
rect 556 581 590 615
rect 556 513 590 543
rect 556 509 590 513
rect 556 467 590 471
rect 556 437 590 467
rect 556 365 590 399
rect 556 293 590 327
rect 556 221 590 255
rect 708 745 710 759
rect 710 745 742 759
rect 708 725 742 745
rect 708 677 710 687
rect 710 677 742 687
rect 708 653 742 677
rect 708 609 710 615
rect 710 609 742 615
rect 708 581 742 609
rect 708 541 710 543
rect 710 541 742 543
rect 708 509 742 541
rect 708 439 742 471
rect 708 437 710 439
rect 710 437 742 439
rect 708 371 742 399
rect 708 365 710 371
rect 710 365 742 371
rect 708 303 742 327
rect 708 293 710 303
rect 710 293 742 303
rect 708 235 742 255
rect 708 221 710 235
rect 710 221 742 235
rect 255 123 289 125
rect 337 123 371 125
rect 431 123 465 125
rect 513 123 547 125
rect 255 91 264 123
rect 264 91 289 123
rect 337 91 371 123
rect 431 91 465 123
rect 513 91 538 123
rect 538 91 547 123
rect 255 19 289 53
rect 337 19 371 53
rect 431 19 465 53
rect 513 19 547 53
<< metal1 >>
rect 243 961 559 980
rect 243 927 255 961
rect 289 927 337 961
rect 371 927 431 961
rect 465 927 513 961
rect 547 927 559 961
rect 243 889 559 927
rect 243 855 255 889
rect 289 855 337 889
rect 371 855 431 889
rect 465 855 513 889
rect 547 855 559 889
rect 243 843 559 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 203 759 255 771
rect 203 725 212 759
rect 246 725 255 759
rect 203 687 255 725
rect 203 653 212 687
rect 246 653 255 687
rect 203 615 255 653
rect 203 581 212 615
rect 246 581 255 615
rect 203 543 255 581
rect 203 509 212 543
rect 246 509 255 543
rect 203 471 255 509
rect 203 459 212 471
rect 246 459 255 471
rect 203 399 255 407
rect 203 395 212 399
rect 246 395 255 399
rect 203 331 255 343
rect 203 267 255 279
rect 203 209 255 215
rect 289 765 341 771
rect 289 701 341 713
rect 289 637 341 649
rect 289 581 298 585
rect 332 581 341 585
rect 289 573 341 581
rect 289 509 298 521
rect 332 509 341 521
rect 289 471 341 509
rect 289 437 298 471
rect 332 437 341 471
rect 289 399 341 437
rect 289 365 298 399
rect 332 365 341 399
rect 289 327 341 365
rect 289 293 298 327
rect 332 293 341 327
rect 289 255 341 293
rect 289 221 298 255
rect 332 221 341 255
rect 289 209 341 221
rect 375 759 427 771
rect 375 725 384 759
rect 418 725 427 759
rect 375 687 427 725
rect 375 653 384 687
rect 418 653 427 687
rect 375 615 427 653
rect 375 581 384 615
rect 418 581 427 615
rect 375 543 427 581
rect 375 509 384 543
rect 418 509 427 543
rect 375 471 427 509
rect 375 459 384 471
rect 418 459 427 471
rect 375 399 427 407
rect 375 395 384 399
rect 418 395 427 399
rect 375 331 427 343
rect 375 267 427 279
rect 375 209 427 215
rect 461 765 513 771
rect 461 701 513 713
rect 461 637 513 649
rect 461 581 470 585
rect 504 581 513 585
rect 461 573 513 581
rect 461 509 470 521
rect 504 509 513 521
rect 461 471 513 509
rect 461 437 470 471
rect 504 437 513 471
rect 461 399 513 437
rect 461 365 470 399
rect 504 365 513 399
rect 461 327 513 365
rect 461 293 470 327
rect 504 293 513 327
rect 461 255 513 293
rect 461 221 470 255
rect 504 221 513 255
rect 461 209 513 221
rect 547 759 599 771
rect 547 725 556 759
rect 590 725 599 759
rect 547 687 599 725
rect 547 653 556 687
rect 590 653 599 687
rect 547 615 599 653
rect 547 581 556 615
rect 590 581 599 615
rect 547 543 599 581
rect 547 509 556 543
rect 590 509 599 543
rect 547 471 599 509
rect 547 459 556 471
rect 590 459 599 471
rect 547 399 599 407
rect 547 395 556 399
rect 590 395 599 399
rect 547 331 599 343
rect 547 267 599 279
rect 547 209 599 215
rect 702 759 761 771
rect 702 725 708 759
rect 742 725 761 759
rect 702 687 761 725
rect 702 653 708 687
rect 742 653 761 687
rect 702 615 761 653
rect 702 581 708 615
rect 742 581 761 615
rect 702 543 761 581
rect 702 509 708 543
rect 742 509 761 543
rect 702 471 761 509
rect 702 437 708 471
rect 742 437 761 471
rect 702 399 761 437
rect 702 365 708 399
rect 742 365 761 399
rect 702 327 761 365
rect 702 293 708 327
rect 742 293 761 327
rect 702 255 761 293
rect 702 221 708 255
rect 742 221 761 255
rect 702 209 761 221
rect 243 125 559 137
rect 243 91 255 125
rect 289 91 337 125
rect 371 91 431 125
rect 465 91 513 125
rect 547 91 559 125
rect 243 53 559 91
rect 243 19 255 53
rect 289 19 337 53
rect 371 19 431 53
rect 465 19 513 53
rect 547 19 559 53
rect 243 0 559 19
<< via1 >>
rect 203 437 212 459
rect 212 437 246 459
rect 246 437 255 459
rect 203 407 255 437
rect 203 365 212 395
rect 212 365 246 395
rect 246 365 255 395
rect 203 343 255 365
rect 203 327 255 331
rect 203 293 212 327
rect 212 293 246 327
rect 246 293 255 327
rect 203 279 255 293
rect 203 255 255 267
rect 203 221 212 255
rect 212 221 246 255
rect 246 221 255 255
rect 203 215 255 221
rect 289 759 341 765
rect 289 725 298 759
rect 298 725 332 759
rect 332 725 341 759
rect 289 713 341 725
rect 289 687 341 701
rect 289 653 298 687
rect 298 653 332 687
rect 332 653 341 687
rect 289 649 341 653
rect 289 615 341 637
rect 289 585 298 615
rect 298 585 332 615
rect 332 585 341 615
rect 289 543 341 573
rect 289 521 298 543
rect 298 521 332 543
rect 332 521 341 543
rect 375 437 384 459
rect 384 437 418 459
rect 418 437 427 459
rect 375 407 427 437
rect 375 365 384 395
rect 384 365 418 395
rect 418 365 427 395
rect 375 343 427 365
rect 375 327 427 331
rect 375 293 384 327
rect 384 293 418 327
rect 418 293 427 327
rect 375 279 427 293
rect 375 255 427 267
rect 375 221 384 255
rect 384 221 418 255
rect 418 221 427 255
rect 375 215 427 221
rect 461 759 513 765
rect 461 725 470 759
rect 470 725 504 759
rect 504 725 513 759
rect 461 713 513 725
rect 461 687 513 701
rect 461 653 470 687
rect 470 653 504 687
rect 504 653 513 687
rect 461 649 513 653
rect 461 615 513 637
rect 461 585 470 615
rect 470 585 504 615
rect 504 585 513 615
rect 461 543 513 573
rect 461 521 470 543
rect 470 521 504 543
rect 504 521 513 543
rect 547 437 556 459
rect 556 437 590 459
rect 590 437 599 459
rect 547 407 599 437
rect 547 365 556 395
rect 556 365 590 395
rect 590 365 599 395
rect 547 343 599 365
rect 547 327 599 331
rect 547 293 556 327
rect 556 293 590 327
rect 590 293 599 327
rect 547 279 599 293
rect 547 255 599 267
rect 547 221 556 255
rect 556 221 590 255
rect 590 221 599 255
rect 547 215 599 221
<< metal2 >>
rect 14 765 788 771
rect 14 713 289 765
rect 341 713 461 765
rect 513 713 788 765
rect 14 701 788 713
rect 14 649 289 701
rect 341 649 461 701
rect 513 649 788 701
rect 14 637 788 649
rect 14 585 289 637
rect 341 585 461 637
rect 513 585 788 637
rect 14 573 788 585
rect 14 521 289 573
rect 341 521 461 573
rect 513 521 788 573
rect 14 515 788 521
rect 14 459 788 465
rect 14 407 203 459
rect 255 407 375 459
rect 427 407 547 459
rect 599 407 788 459
rect 14 395 788 407
rect 14 343 203 395
rect 255 343 375 395
rect 427 343 547 395
rect 599 343 788 395
rect 14 331 788 343
rect 14 279 203 331
rect 255 279 375 331
rect 427 279 547 331
rect 599 279 788 331
rect 14 267 788 279
rect 14 215 203 267
rect 255 215 375 267
rect 427 215 547 267
rect 599 215 788 267
rect 14 209 788 215
<< labels >>
flabel metal1 s 301 878 511 928 0 FreeSans 200 0 0 0 GATE
port 4 nsew
flabel metal1 s 301 42 511 92 0 FreeSans 200 0 0 0 GATE
port 4 nsew
flabel metal1 s 41 466 100 496 0 FreeSans 200 90 0 0 SUBSTRATE
port 3 nsew
flabel metal1 s 702 469 761 499 0 FreeSans 200 90 0 0 SUBSTRATE
port 3 nsew
flabel comment s 229 490 229 490 0 FreeSans 300 0 0 0 S
flabel comment s 315 490 315 490 0 FreeSans 300 0 0 0 S
flabel comment s 401 490 401 490 0 FreeSans 300 0 0 0 S
flabel comment s 487 490 487 490 0 FreeSans 300 0 0 0 S
flabel comment s 229 490 229 490 0 FreeSans 300 0 0 0 S
flabel comment s 315 490 315 490 0 FreeSans 300 0 0 0 D
flabel comment s 401 490 401 490 0 FreeSans 300 0 0 0 S
flabel comment s 487 490 487 490 0 FreeSans 300 0 0 0 D
flabel comment s 573 490 573 490 0 FreeSans 300 0 0 0 S
flabel comment s 182 496 182 496 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 613 488 613 488 0 FreeSans 180 90 0 0 dummy_poly
flabel metal2 s 14 280 35 408 7 FreeSans 300 180 0 0 SOURCE
port 5 nsew
flabel metal2 s 14 589 35 717 7 FreeSans 300 180 0 0 DRAIN
port 6 nsew
<< properties >>
string GDS_END 6687678
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6670436
<< end >>
