magic
tech sky130B
magscale 1 2
timestamp 1686671242
<< nwell >>
rect -36 679 1268 1471
<< locali >>
rect 0 1397 1232 1431
rect 64 674 98 740
rect 613 690 647 724
rect 0 -17 1232 17
use sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_14  sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_14_0
timestamp 1686671242
transform 1 0 0 0 1 0
box -36 -17 1268 1471
<< labels >>
rlabel locali s 630 707 630 707 4 Z
rlabel locali s 81 707 81 707 4 A
rlabel locali s 616 0 616 0 4 gnd
rlabel locali s 616 1414 616 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1232 1414
string GDS_END 323046
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 322214
<< end >>
