magic
tech sky130B
magscale 1 2
timestamp 1686671242
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_0
timestamp 1686671242
transform -1 0 -80 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_1
timestamp 1686671242
transform 1 0 117 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 15438276
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 15437286
<< end >>
