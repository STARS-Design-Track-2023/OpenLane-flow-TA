magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< locali >>
rect 356 1137 390 1153
rect 10340 1137 10374 1153
rect 20324 1137 20358 1153
rect 30308 1137 30342 1153
rect 0 1103 356 1137
rect 390 1103 10340 1137
rect 10374 1103 20324 1137
rect 20358 1103 30308 1137
rect 30342 1103 30698 1137
rect 356 1087 390 1103
rect 10340 1087 10374 1103
rect 20324 1087 20358 1103
rect 30308 1087 30342 1103
rect 212 535 246 551
rect 557 524 591 558
rect 10196 535 10230 551
rect 212 485 246 501
rect 10541 524 10575 558
rect 20180 535 20214 551
rect 10196 485 10230 501
rect 20525 524 20559 558
rect 30164 535 30198 551
rect 20180 485 20214 501
rect 30509 524 30543 558
rect 30164 485 30198 501
rect -17 287 17 303
rect 9967 287 10001 303
rect 19951 287 19985 303
rect 29935 287 29969 303
rect 17 253 129 287
rect 10001 253 10113 287
rect 19985 253 20097 287
rect 29969 253 30081 287
rect -17 237 17 253
rect 9967 237 10001 253
rect 19951 237 19985 253
rect 29935 237 29969 253
rect 356 17 390 33
rect 10340 17 10374 33
rect 20324 17 20358 33
rect 30308 17 30342 33
rect 0 -17 356 17
rect 390 -17 10340 17
rect 10374 -17 20324 17
rect 20358 -17 30308 17
rect 30342 -17 30698 17
rect 356 -33 390 -17
rect 10340 -33 10374 -17
rect 20324 -33 20358 -17
rect 30308 -33 30342 -17
<< viali >>
rect 356 1103 390 1137
rect 10340 1103 10374 1137
rect 20324 1103 20358 1137
rect 30308 1103 30342 1137
rect 212 501 246 535
rect 10196 501 10230 535
rect 20180 501 20214 535
rect 30164 501 30198 535
rect -17 253 17 287
rect 9967 253 10001 287
rect 19951 253 19985 287
rect 29935 253 29969 287
rect 356 -17 390 17
rect 10340 -17 10374 17
rect 20324 -17 20358 17
rect 30308 -17 30342 17
<< metal1 >>
rect 341 1094 347 1146
rect 399 1094 405 1146
rect 10325 1094 10331 1146
rect 10383 1094 10389 1146
rect 20309 1094 20315 1146
rect 20367 1094 20373 1146
rect 30293 1094 30299 1146
rect 30351 1094 30357 1146
rect 197 492 203 544
rect 255 492 261 544
rect 10181 492 10187 544
rect 10239 492 10245 544
rect 20165 492 20171 544
rect 20223 492 20229 544
rect 30149 492 30155 544
rect 30207 492 30213 544
rect -32 244 -26 296
rect 26 244 32 296
rect 9952 244 9958 296
rect 10010 244 10016 296
rect 19936 244 19942 296
rect 19994 244 20000 296
rect 29920 244 29926 296
rect 29978 244 29984 296
rect 341 -26 347 26
rect 399 -26 405 26
rect 10325 -26 10331 26
rect 10383 -26 10389 26
rect 20309 -26 20315 26
rect 20367 -26 20373 26
rect 30293 -26 30299 26
rect 30351 -26 30357 26
<< via1 >>
rect 347 1137 399 1146
rect 347 1103 356 1137
rect 356 1103 390 1137
rect 390 1103 399 1137
rect 347 1094 399 1103
rect 10331 1137 10383 1146
rect 10331 1103 10340 1137
rect 10340 1103 10374 1137
rect 10374 1103 10383 1137
rect 10331 1094 10383 1103
rect 20315 1137 20367 1146
rect 20315 1103 20324 1137
rect 20324 1103 20358 1137
rect 20358 1103 20367 1137
rect 20315 1094 20367 1103
rect 30299 1137 30351 1146
rect 30299 1103 30308 1137
rect 30308 1103 30342 1137
rect 30342 1103 30351 1137
rect 30299 1094 30351 1103
rect 203 535 255 544
rect 203 501 212 535
rect 212 501 246 535
rect 246 501 255 535
rect 203 492 255 501
rect 10187 535 10239 544
rect 10187 501 10196 535
rect 10196 501 10230 535
rect 10230 501 10239 535
rect 10187 492 10239 501
rect 20171 535 20223 544
rect 20171 501 20180 535
rect 20180 501 20214 535
rect 20214 501 20223 535
rect 20171 492 20223 501
rect 30155 535 30207 544
rect 30155 501 30164 535
rect 30164 501 30198 535
rect 30198 501 30207 535
rect 30155 492 30207 501
rect -26 287 26 296
rect -26 253 -17 287
rect -17 253 17 287
rect 17 253 26 287
rect -26 244 26 253
rect 9958 287 10010 296
rect 9958 253 9967 287
rect 9967 253 10001 287
rect 10001 253 10010 287
rect 9958 244 10010 253
rect 19942 287 19994 296
rect 19942 253 19951 287
rect 19951 253 19985 287
rect 19985 253 19994 287
rect 19942 244 19994 253
rect 29926 287 29978 296
rect 29926 253 29935 287
rect 29935 253 29969 287
rect 29969 253 29978 287
rect 29926 244 29978 253
rect 347 17 399 26
rect 347 -17 356 17
rect 356 -17 390 17
rect 390 -17 399 17
rect 347 -26 399 -17
rect 10331 17 10383 26
rect 10331 -17 10340 17
rect 10340 -17 10374 17
rect 10374 -17 10383 17
rect 10331 -26 10383 -17
rect 20315 17 20367 26
rect 20315 -17 20324 17
rect 20324 -17 20358 17
rect 20358 -17 20367 17
rect 20315 -26 20367 -17
rect 30299 17 30351 26
rect 30299 -17 30308 17
rect 30308 -17 30342 17
rect 30342 -17 30351 17
rect 30299 -26 30351 -17
<< metal2 >>
rect 345 1148 401 1157
rect 345 1083 401 1092
rect 10329 1148 10385 1157
rect 10329 1083 10385 1092
rect 20313 1148 20369 1157
rect 20313 1083 20369 1092
rect 30297 1148 30353 1157
rect 30297 1083 30353 1092
rect 201 546 257 555
rect 201 481 257 490
rect 10185 546 10241 555
rect 10185 481 10241 490
rect 20169 546 20225 555
rect 20169 481 20225 490
rect 30153 546 30209 555
rect 30153 481 30209 490
rect -26 296 26 302
rect -26 238 26 244
rect 9958 296 10010 302
rect 9958 238 10010 244
rect 19942 296 19994 302
rect 19942 238 19994 244
rect 29926 296 29978 302
rect 29926 238 29978 244
rect 345 28 401 37
rect 345 -37 401 -28
rect 10329 28 10385 37
rect 10329 -37 10385 -28
rect 20313 28 20369 37
rect 20313 -37 20369 -28
rect 30297 28 30353 37
rect 30297 -37 30353 -28
<< via2 >>
rect 345 1146 401 1148
rect 345 1094 347 1146
rect 347 1094 399 1146
rect 399 1094 401 1146
rect 345 1092 401 1094
rect 10329 1146 10385 1148
rect 10329 1094 10331 1146
rect 10331 1094 10383 1146
rect 10383 1094 10385 1146
rect 10329 1092 10385 1094
rect 20313 1146 20369 1148
rect 20313 1094 20315 1146
rect 20315 1094 20367 1146
rect 20367 1094 20369 1146
rect 20313 1092 20369 1094
rect 30297 1146 30353 1148
rect 30297 1094 30299 1146
rect 30299 1094 30351 1146
rect 30351 1094 30353 1146
rect 30297 1092 30353 1094
rect 201 544 257 546
rect 201 492 203 544
rect 203 492 255 544
rect 255 492 257 544
rect 201 490 257 492
rect 10185 544 10241 546
rect 10185 492 10187 544
rect 10187 492 10239 544
rect 10239 492 10241 544
rect 10185 490 10241 492
rect 20169 544 20225 546
rect 20169 492 20171 544
rect 20171 492 20223 544
rect 20223 492 20225 544
rect 20169 490 20225 492
rect 30153 544 30209 546
rect 30153 492 30155 544
rect 30155 492 30207 544
rect 30207 492 30209 544
rect 30153 490 30209 492
rect 345 26 401 28
rect 345 -26 347 26
rect 347 -26 399 26
rect 399 -26 401 26
rect 345 -28 401 -26
rect 10329 26 10385 28
rect 10329 -26 10331 26
rect 10331 -26 10383 26
rect 10383 -26 10385 26
rect 10329 -28 10385 -26
rect 20313 26 20369 28
rect 20313 -26 20315 26
rect 20315 -26 20367 26
rect 20367 -26 20369 26
rect 20313 -28 20369 -26
rect 30297 26 30353 28
rect 30297 -26 30299 26
rect 30299 -26 30351 26
rect 30351 -26 30353 26
rect 30297 -28 30353 -26
<< metal3 >>
rect 324 1148 422 1169
rect 324 1092 345 1148
rect 401 1092 422 1148
rect 324 1071 422 1092
rect 10308 1148 10406 1169
rect 10308 1092 10329 1148
rect 10385 1092 10406 1148
rect 10308 1071 10406 1092
rect 20292 1148 20390 1169
rect 20292 1092 20313 1148
rect 20369 1092 20390 1148
rect 20292 1071 20390 1092
rect 30276 1148 30374 1169
rect 30276 1092 30297 1148
rect 30353 1092 30374 1148
rect 30276 1071 30374 1092
rect 196 548 262 551
rect 10180 548 10246 551
rect 20164 548 20230 551
rect 30148 548 30214 551
rect 0 546 39936 548
rect 0 490 201 546
rect 257 490 10185 546
rect 10241 490 20169 546
rect 20225 490 30153 546
rect 30209 490 39936 546
rect 0 488 39936 490
rect 196 485 262 488
rect 10180 485 10246 488
rect 20164 485 20230 488
rect 30148 485 30214 488
rect 324 28 422 49
rect 324 -28 345 28
rect 401 -28 422 28
rect 324 -49 422 -28
rect 10308 28 10406 49
rect 10308 -28 10329 28
rect 10385 -28 10406 28
rect 10308 -49 10406 -28
rect 20292 28 20390 49
rect 20292 -28 20313 28
rect 20369 -28 20390 28
rect 20292 -49 20390 -28
rect 30276 28 30374 49
rect 30276 -28 30297 28
rect 30353 -28 30374 28
rect 30276 -49 30374 -28
use contact_7  contact_7_0
timestamp 1683767628
transform 1 0 30296 0 1 1087
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1683767628
transform 1 0 30296 0 1 -33
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1683767628
transform 1 0 30152 0 1 485
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1683767628
transform 1 0 29923 0 1 237
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1683767628
transform 1 0 20312 0 1 1087
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1683767628
transform 1 0 20312 0 1 -33
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1683767628
transform 1 0 20168 0 1 485
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1683767628
transform 1 0 19939 0 1 237
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1683767628
transform 1 0 10328 0 1 1087
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1683767628
transform 1 0 10328 0 1 -33
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1683767628
transform 1 0 10184 0 1 485
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1683767628
transform 1 0 9955 0 1 237
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1683767628
transform 1 0 344 0 1 1087
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1683767628
transform 1 0 344 0 1 -33
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1683767628
transform 1 0 200 0 1 485
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1683767628
transform 1 0 -29 0 1 237
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1683767628
transform 1 0 30293 0 1 1088
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1683767628
transform 1 0 30293 0 1 -32
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1683767628
transform 1 0 30149 0 1 486
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1683767628
transform 1 0 29920 0 1 238
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1683767628
transform 1 0 20309 0 1 1088
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1683767628
transform 1 0 20309 0 1 -32
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1683767628
transform 1 0 20165 0 1 486
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1683767628
transform 1 0 19936 0 1 238
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1683767628
transform 1 0 10325 0 1 1088
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1683767628
transform 1 0 10325 0 1 -32
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1683767628
transform 1 0 10181 0 1 486
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1683767628
transform 1 0 9952 0 1 238
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1683767628
transform 1 0 341 0 1 1088
box 0 0 1 1
use contact_8  contact_8_13
timestamp 1683767628
transform 1 0 341 0 1 -32
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1683767628
transform 1 0 197 0 1 486
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1683767628
transform 1 0 -32 0 1 238
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1683767628
transform 1 0 30292 0 1 1083
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1683767628
transform 1 0 30292 0 1 -37
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1683767628
transform 1 0 30148 0 1 481
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1683767628
transform 1 0 20308 0 1 1083
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1683767628
transform 1 0 20308 0 1 -37
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1683767628
transform 1 0 20164 0 1 481
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1683767628
transform 1 0 10324 0 1 1083
box 0 0 1 1
use contact_9  contact_9_7
timestamp 1683767628
transform 1 0 10324 0 1 -37
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1683767628
transform 1 0 10180 0 1 481
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1683767628
transform 1 0 340 0 1 1083
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1683767628
transform 1 0 340 0 1 -37
box 0 0 1 1
use contact_9  contact_9_11
timestamp 1683767628
transform 1 0 196 0 1 481
box 0 0 1 1
use pand2  pand2_0
timestamp 1683767628
transform 1 0 29952 0 1 0
box -36 -17 782 1177
use pand2  pand2_1
timestamp 1683767628
transform 1 0 19968 0 1 0
box -36 -17 782 1177
use pand2  pand2_2
timestamp 1683767628
transform 1 0 9984 0 1 0
box -36 -17 782 1177
use pand2  pand2_3
timestamp 1683767628
transform 1 0 0 0 1 0
box -36 -17 782 1177
<< labels >>
rlabel locali s 10558 541 10558 541 4 wmask_out_1
port 7 nsew
rlabel locali s 20542 541 20542 541 4 wmask_out_2
port 8 nsew
rlabel locali s 30526 541 30526 541 4 wmask_out_3
port 9 nsew
rlabel locali s 574 541 574 541 4 wmask_out_0
port 6 nsew
rlabel metal2 s 19968 270 19968 270 4 wmask_in_2
port 3 nsew
rlabel metal2 s 9984 270 9984 270 4 wmask_in_1
port 2 nsew
rlabel metal2 s 0 270 0 270 4 wmask_in_0
port 1 nsew
rlabel metal2 s 29952 270 29952 270 4 wmask_in_3
port 4 nsew
rlabel metal3 s 20341 1120 20341 1120 4 vdd
port 10 nsew
rlabel metal3 s 373 1120 373 1120 4 vdd
port 10 nsew
rlabel metal3 s 10357 1120 10357 1120 4 vdd
port 10 nsew
rlabel metal3 s 30325 1120 30325 1120 4 vdd
port 10 nsew
rlabel metal3 s 30325 0 30325 0 4 gnd
port 11 nsew
rlabel metal3 s 10357 0 10357 0 4 gnd
port 11 nsew
rlabel metal3 s 373 0 373 0 4 gnd
port 11 nsew
rlabel metal3 s 20341 0 20341 0 4 gnd
port 11 nsew
rlabel metal3 s 19968 518 19968 518 4 en
port 5 nsew
<< properties >>
string FIXED_BBOX 30292 -37 30358 0
string GDS_END 3513744
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 3507692
<< end >>
